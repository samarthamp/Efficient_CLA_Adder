magic
tech scmos
timestamp 1731176518
<< nwell >>
rect -39 21 -15 53
rect 0 0 60 52
rect -39 -58 -15 -26
<< ntransistor >>
rect -28 4 -26 14
rect -28 -19 -26 -9
rect 11 -44 13 -14
rect 21 -44 23 -14
rect 37 -44 39 -14
rect 47 -44 49 -14
<< ptransistor >>
rect -28 27 -26 47
rect 11 6 13 46
rect 21 6 23 46
rect 37 6 39 46
rect 47 6 49 46
rect -28 -52 -26 -32
<< ndiffusion >>
rect -33 8 -28 14
rect -29 4 -28 8
rect -26 10 -25 14
rect -26 4 -21 10
rect -29 -13 -28 -9
rect -33 -19 -28 -13
rect -26 -15 -21 -9
rect -26 -19 -25 -15
rect 6 -40 11 -14
rect 10 -44 11 -40
rect 13 -44 21 -14
rect 23 -18 28 -14
rect 32 -18 37 -14
rect 23 -44 37 -18
rect 39 -44 47 -14
rect 49 -40 54 -14
rect 49 -44 50 -40
<< pdiffusion >>
rect -29 43 -28 47
rect -33 27 -28 43
rect -26 31 -21 47
rect -26 27 -25 31
rect 10 42 11 46
rect 6 6 11 42
rect 13 10 21 46
rect 13 6 15 10
rect 19 6 21 10
rect 23 42 24 46
rect 23 6 28 42
rect 36 42 37 46
rect 32 10 37 42
rect 36 6 37 10
rect 39 10 47 46
rect 39 6 41 10
rect 45 6 47 10
rect 49 42 50 46
rect 49 6 54 42
rect -33 -48 -28 -32
rect -29 -52 -28 -48
rect -26 -36 -25 -32
rect -26 -52 -21 -36
<< ndcontact >>
rect -33 4 -29 8
rect -25 10 -21 14
rect -33 -13 -29 -9
rect -25 -19 -21 -15
rect 6 -44 10 -40
rect 28 -18 32 -14
rect 50 -44 54 -40
<< pdcontact >>
rect -33 43 -29 47
rect -25 27 -21 31
rect 6 42 10 46
rect 15 6 19 10
rect 24 42 28 46
rect 32 42 36 46
rect 32 6 36 10
rect 41 6 45 10
rect 50 42 54 46
rect -33 -52 -29 -48
rect -25 -36 -21 -32
<< polysilicon >>
rect -28 47 -26 51
rect 11 46 13 49
rect 21 46 23 49
rect 37 46 39 59
rect 47 46 49 49
rect -28 14 -26 27
rect -28 0 -26 4
rect 11 -1 13 6
rect -28 -9 -26 -5
rect 11 -14 13 -6
rect 21 -8 23 6
rect 21 -14 23 -13
rect 37 -14 39 6
rect 47 -14 49 6
rect -28 -32 -26 -19
rect 11 -47 13 -44
rect 21 -47 23 -44
rect 37 -47 39 -44
rect -28 -56 -26 -52
rect 47 -54 49 -44
<< polycontact >>
rect -32 15 -28 19
rect -32 -24 -28 -20
<< metal1 >>
rect -45 54 28 57
rect -45 -59 -42 54
rect -33 47 -29 54
rect 6 46 10 54
rect 24 46 28 54
rect 32 53 54 56
rect 32 46 36 53
rect 50 46 54 53
rect -25 20 -21 27
rect -34 15 -32 19
rect -25 14 -21 15
rect -33 -1 -29 4
rect 16 -1 19 6
rect 32 -1 36 6
rect -33 -4 -7 -1
rect -33 -9 -29 -4
rect -25 -20 -21 -19
rect -34 -24 -32 -20
rect -25 -32 -21 -25
rect -10 -48 -7 -4
rect 16 -4 36 -1
rect 41 -8 45 6
rect 28 -11 60 -8
rect 28 -14 32 -11
rect 6 -48 10 -44
rect 50 -48 54 -44
rect -10 -51 54 -48
rect -33 -59 -29 -52
rect -45 -62 -29 -59
<< m2contact >>
rect -39 14 -34 19
rect -25 15 -20 20
rect -39 -24 -34 -19
rect -25 -25 -20 -20
<< pm12contact >>
rect 34 59 39 64
rect 8 -6 13 -1
rect 18 -13 23 -8
rect 44 -59 49 -54
<< metal2 >>
rect -4 59 34 64
rect -4 20 -1 59
rect -20 15 -1 20
rect -39 -1 -36 14
rect -39 -4 8 -1
rect -39 -13 18 -10
rect -39 -19 -36 -13
rect -20 -25 -1 -20
rect -4 -54 -1 -25
rect -4 -59 44 -54
<< labels >>
rlabel metal1 -32 1 -30 3 1 gnd
rlabel metal1 -32 54 -30 56 5 vdd
rlabel m2contact -38 -23 -36 -21 1 b
rlabel m2contact -38 16 -36 18 1 a
rlabel metal2 -14 16 -12 18 1 a_bar
rlabel metal2 -15 -23 -13 -22 1 b_bar
rlabel metal1 55 -10 58 -9 7 out
<< end >>
