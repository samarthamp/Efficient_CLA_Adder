magic
tech scmos
timestamp 1731162172
<< nwell >>
rect 0 -20 34 32
<< ntransistor >>
rect 11 -43 13 -33
rect 21 -43 23 -33
<< ptransistor >>
rect 11 -14 13 26
rect 21 -14 23 26
<< ndiffusion >>
rect 6 -39 11 -33
rect 10 -43 11 -39
rect 13 -37 15 -33
rect 19 -37 21 -33
rect 13 -43 21 -37
rect 23 -39 28 -33
rect 23 -43 24 -39
<< pdiffusion >>
rect 10 22 11 26
rect 6 -14 11 22
rect 13 -14 21 26
rect 23 -10 28 26
rect 23 -14 24 -10
<< ndcontact >>
rect 6 -43 10 -39
rect 15 -37 19 -33
rect 24 -43 28 -39
<< pdcontact >>
rect 6 22 10 26
rect 24 -14 28 -10
<< polysilicon >>
rect 11 26 13 29
rect 21 26 23 29
rect 11 -33 13 -14
rect 21 -33 23 -14
rect 11 -46 13 -43
rect 21 -46 23 -43
<< polycontact >>
rect 7 -32 11 -28
rect 17 -25 21 -21
<< metal1 >>
rect 6 26 10 36
rect 0 -25 17 -21
rect 24 -28 28 -14
rect 0 -32 7 -28
rect 15 -32 34 -28
rect 15 -33 19 -32
rect 6 -47 10 -43
rect 24 -47 28 -43
rect 6 -50 28 -47
<< labels >>
rlabel metal1 3 -31 4 -30 3 a
rlabel metal1 4 -24 6 -22 3 b
rlabel metal1 30 -31 32 -29 7 out
rlabel metal1 7 33 8 35 5 vdd
rlabel metal1 16 -49 17 -48 1 gnd
<< end >>
