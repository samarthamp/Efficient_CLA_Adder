magic
tech scmos
timestamp 1731503625
<< nwell >>
rect 318 -146 370 -82
rect 378 -119 402 -87
rect 409 -119 433 -87
rect 441 -146 493 -82
rect 318 -162 350 -146
rect 318 -192 350 -168
rect 357 -188 381 -156
rect 430 -188 454 -156
rect 461 -162 493 -146
rect 461 -192 493 -168
rect 189 -256 221 -232
rect 258 -235 290 -211
rect 231 -263 295 -243
rect 141 -295 165 -263
rect 185 -295 209 -263
rect 215 -295 295 -263
rect 337 -275 369 -241
rect 437 -275 489 -241
rect 31 -326 63 -302
rect 331 -318 365 -286
rect 26 -354 90 -334
rect 100 -347 132 -323
rect 372 -337 424 -285
rect 569 -290 649 -258
rect 655 -290 679 -258
rect 699 -290 723 -258
rect 748 -279 780 -255
rect 569 -310 633 -290
rect 26 -386 106 -354
rect 112 -386 136 -354
rect 465 -359 489 -327
rect 574 -342 606 -318
rect 643 -321 675 -297
rect 743 -307 807 -287
rect 817 -300 849 -276
rect 743 -339 823 -307
rect 829 -339 853 -307
rect 873 -339 897 -307
rect 196 -404 228 -380
rect 251 -404 283 -361
rect 446 -414 489 -382
rect -113 -463 -33 -431
rect -27 -463 -3 -431
rect -113 -483 -49 -463
rect -108 -515 -76 -491
rect -39 -494 -7 -470
rect 42 -486 76 -434
rect 196 -469 228 -445
rect 251 -469 283 -426
rect 338 -447 362 -415
rect 550 -422 602 -370
rect 616 -382 648 -348
rect 616 -426 668 -391
rect -108 -545 -76 -521
rect -113 -573 -49 -553
rect -39 -566 -7 -542
rect 116 -546 168 -494
rect 181 -528 233 -494
rect 319 -502 362 -470
rect 398 -507 422 -475
rect 570 -483 602 -433
rect 616 -467 648 -433
rect 708 -466 742 -434
rect 786 -463 810 -431
rect 816 -463 896 -431
rect 440 -519 472 -485
rect 551 -526 603 -492
rect 616 -526 668 -474
rect 790 -494 822 -470
rect 832 -483 896 -463
rect 859 -515 891 -491
rect -113 -605 -33 -573
rect -27 -605 -3 -573
rect 42 -586 76 -554
rect 136 -587 168 -553
rect 182 -587 214 -537
rect 489 -585 532 -553
rect 116 -646 168 -594
rect 205 -645 237 -602
rect 260 -650 292 -602
rect 315 -650 347 -607
rect 398 -640 432 -588
rect 627 -599 659 -575
rect 708 -586 742 -534
rect 790 -566 822 -542
rect 859 -545 891 -521
rect 832 -573 896 -553
rect 441 -639 491 -607
rect 508 -640 532 -608
rect 565 -652 589 -620
rect 622 -627 686 -607
rect 696 -620 728 -596
rect 786 -605 810 -573
rect 816 -605 896 -573
rect 398 -705 450 -653
rect 457 -685 491 -653
rect 498 -705 550 -653
rect 622 -659 702 -627
rect 708 -659 732 -627
rect 752 -659 776 -627
rect 565 -707 608 -675
rect 177 -751 201 -719
rect 221 -751 245 -719
rect 251 -751 331 -719
rect 225 -782 257 -758
rect 267 -771 331 -751
rect 337 -779 389 -745
rect 457 -779 489 -745
rect 294 -803 326 -779
rect 350 -846 382 -822
rect 350 -868 382 -852
rect 389 -858 413 -826
rect 461 -858 485 -826
rect 492 -846 524 -822
rect 492 -868 524 -852
rect 350 -932 402 -868
rect 410 -927 434 -895
rect 440 -927 464 -895
rect 472 -932 524 -868
<< ntransistor >>
rect 293 -95 303 -93
rect 508 -95 518 -93
rect 293 -121 303 -119
rect 508 -121 518 -119
rect 389 -135 391 -125
rect 420 -135 422 -125
rect 292 -151 312 -149
rect 499 -151 519 -149
rect 292 -161 312 -159
rect 499 -161 519 -159
rect 292 -181 312 -179
rect 499 -181 519 -179
rect 292 -191 312 -189
rect 499 -191 519 -189
rect 368 -204 370 -194
rect 441 -204 443 -194
rect 242 -224 252 -222
rect 580 -243 582 -233
rect 173 -245 183 -243
rect 383 -254 403 -252
rect 414 -254 424 -252
rect 383 -264 403 -262
rect 414 -264 424 -262
rect 606 -243 608 -233
rect 636 -252 638 -232
rect 646 -252 648 -232
rect 666 -252 668 -232
rect 676 -252 678 -232
rect 710 -252 712 -242
rect 152 -311 154 -301
rect 69 -315 79 -313
rect 186 -321 188 -301
rect 196 -321 198 -301
rect 216 -321 218 -301
rect 226 -321 228 -301
rect 138 -336 148 -334
rect 256 -320 258 -310
rect 282 -320 284 -310
rect 786 -268 796 -266
rect 855 -289 865 -287
rect 681 -310 691 -308
rect 342 -352 344 -332
rect 352 -352 354 -332
rect 383 -353 385 -343
rect 612 -331 622 -329
rect 401 -360 403 -350
rect 411 -360 413 -350
rect 662 -361 682 -359
rect 289 -374 299 -372
rect 476 -376 478 -366
rect 754 -364 756 -354
rect 662 -371 682 -369
rect -102 -416 -100 -406
rect -76 -416 -74 -406
rect -46 -425 -44 -405
rect -36 -425 -34 -405
rect -16 -425 -14 -405
rect -6 -425 -4 -405
rect 37 -411 39 -401
rect 63 -411 65 -401
rect 534 -383 544 -381
rect 780 -364 782 -354
rect 810 -365 812 -345
rect 820 -365 822 -345
rect 840 -365 842 -345
rect 850 -365 852 -345
rect 884 -355 886 -345
rect 93 -412 95 -392
rect 103 -412 105 -392
rect 123 -412 125 -392
rect 133 -412 135 -392
rect 235 -393 245 -391
rect 289 -393 299 -391
rect 527 -401 537 -399
rect 681 -405 691 -403
rect 527 -411 537 -409
rect 681 -415 691 -413
rect 289 -439 299 -437
rect 457 -430 459 -420
rect 476 -430 478 -420
rect 787 -425 789 -405
rect 797 -425 799 -405
rect 817 -425 819 -405
rect 827 -425 829 -405
rect 857 -416 859 -406
rect 883 -416 885 -406
rect 554 -446 564 -444
rect 662 -446 682 -444
rect 235 -458 245 -456
rect 289 -458 299 -456
rect 349 -464 351 -454
rect 662 -456 682 -454
rect 536 -462 556 -460
rect 536 -472 556 -470
rect -1 -483 9 -481
rect -70 -504 -60 -502
rect 53 -509 55 -499
rect 63 -509 65 -499
rect 93 -507 103 -505
rect 246 -507 256 -505
rect 674 -487 684 -485
rect 486 -498 506 -496
rect 93 -517 103 -515
rect 246 -517 256 -515
rect -70 -534 -60 -532
rect 53 -540 55 -520
rect 63 -540 65 -520
rect 330 -518 332 -508
rect 349 -518 351 -508
rect 719 -500 721 -480
rect 729 -500 731 -480
rect 774 -483 784 -481
rect 528 -505 538 -503
rect 681 -505 691 -503
rect 843 -504 853 -502
rect 486 -508 506 -506
rect 409 -523 411 -513
rect 528 -515 538 -513
rect 681 -515 691 -513
rect 719 -521 721 -511
rect 729 -521 731 -511
rect 100 -535 110 -533
rect -1 -555 9 -553
rect 500 -547 502 -537
rect 519 -547 521 -537
rect 843 -534 853 -532
rect 228 -550 248 -548
rect 228 -560 248 -558
rect 102 -566 122 -564
rect 102 -576 122 -574
rect 220 -576 230 -574
rect 409 -575 411 -565
rect 419 -575 421 -565
rect 452 -593 454 -573
rect 462 -593 464 -573
rect 774 -555 784 -553
rect 665 -588 675 -586
rect -102 -630 -100 -620
rect -76 -630 -74 -620
rect 93 -607 103 -605
rect -46 -631 -44 -611
rect -36 -631 -34 -611
rect -16 -631 -14 -611
rect -6 -631 -4 -611
rect 189 -615 199 -613
rect 243 -615 253 -613
rect 93 -617 103 -615
rect 353 -620 363 -618
rect 100 -635 110 -633
rect 189 -634 199 -632
rect 478 -601 480 -591
rect 519 -601 521 -591
rect 734 -609 744 -607
rect 299 -639 309 -637
rect 353 -639 363 -637
rect 787 -631 789 -611
rect 797 -631 799 -611
rect 817 -631 819 -611
rect 827 -631 829 -611
rect 857 -630 859 -620
rect 883 -630 885 -620
rect 188 -713 190 -703
rect 222 -713 224 -693
rect 232 -713 234 -693
rect 252 -713 254 -693
rect 262 -713 264 -693
rect 292 -704 294 -694
rect 318 -704 320 -694
rect 576 -669 578 -659
rect 409 -728 411 -718
rect 419 -728 421 -718
rect 437 -721 439 -711
rect 468 -719 470 -699
rect 478 -719 480 -699
rect 633 -684 635 -674
rect 509 -728 511 -718
rect 519 -728 521 -718
rect 537 -721 539 -711
rect 659 -684 661 -674
rect 689 -685 691 -665
rect 699 -685 701 -665
rect 719 -685 721 -665
rect 729 -685 731 -665
rect 763 -675 765 -665
rect 576 -723 578 -713
rect 595 -723 597 -713
rect 402 -758 412 -756
rect 423 -758 443 -756
rect 402 -768 412 -766
rect 423 -768 443 -766
rect 209 -771 219 -769
rect 278 -792 288 -790
rect 400 -820 402 -810
rect 472 -820 474 -810
rect 324 -825 344 -823
rect 530 -825 550 -823
rect 324 -835 344 -833
rect 530 -835 550 -833
rect 324 -855 344 -853
rect 530 -855 550 -853
rect 324 -865 344 -863
rect 530 -865 550 -863
rect 421 -889 423 -879
rect 451 -889 453 -879
rect 325 -895 335 -893
rect 539 -895 549 -893
rect 325 -921 335 -919
rect 539 -921 549 -919
<< ptransistor >>
rect 324 -95 364 -93
rect 324 -105 364 -103
rect 389 -113 391 -93
rect 420 -113 422 -93
rect 447 -95 487 -93
rect 447 -105 487 -103
rect 324 -121 364 -119
rect 447 -121 487 -119
rect 324 -131 364 -129
rect 447 -131 487 -129
rect 324 -151 344 -149
rect 467 -151 487 -149
rect 324 -181 344 -179
rect 368 -182 370 -162
rect 441 -182 443 -162
rect 467 -181 487 -179
rect 264 -224 284 -222
rect 195 -245 215 -243
rect 152 -289 154 -269
rect 196 -289 198 -269
rect 226 -289 228 -269
rect 246 -289 248 -249
rect 256 -289 258 -249
rect 272 -289 274 -249
rect 282 -289 284 -249
rect 343 -254 363 -252
rect 443 -254 483 -252
rect 343 -264 363 -262
rect 443 -264 483 -262
rect 37 -315 57 -313
rect 106 -336 126 -334
rect 37 -380 39 -340
rect 47 -380 49 -340
rect 63 -380 65 -340
rect 73 -380 75 -340
rect 342 -312 344 -292
rect 352 -312 354 -292
rect 383 -331 385 -311
rect 401 -331 403 -291
rect 411 -331 413 -291
rect 580 -304 582 -264
rect 590 -304 592 -264
rect 606 -304 608 -264
rect 616 -304 618 -264
rect 636 -284 638 -264
rect 666 -284 668 -264
rect 710 -284 712 -264
rect 754 -268 774 -266
rect 823 -289 843 -287
rect 649 -310 669 -308
rect 580 -331 600 -329
rect 476 -353 478 -333
rect 754 -333 756 -293
rect 764 -333 766 -293
rect 780 -333 782 -293
rect 790 -333 792 -293
rect 810 -333 812 -313
rect 840 -333 842 -313
rect 884 -333 886 -313
rect 93 -380 95 -360
rect 123 -380 125 -360
rect 622 -361 642 -359
rect 257 -374 277 -372
rect 622 -371 642 -369
rect 556 -383 576 -381
rect 202 -393 222 -391
rect 257 -393 277 -391
rect 457 -408 459 -388
rect 476 -408 478 -388
rect 556 -401 596 -399
rect 622 -405 662 -403
rect 556 -411 596 -409
rect 622 -415 662 -413
rect -102 -477 -100 -437
rect -92 -477 -90 -437
rect -76 -477 -74 -437
rect -66 -477 -64 -437
rect -46 -457 -44 -437
rect -16 -457 -14 -437
rect 257 -439 277 -437
rect 53 -480 55 -440
rect 63 -480 65 -440
rect 349 -441 351 -421
rect 576 -446 596 -444
rect 622 -446 642 -444
rect 202 -458 222 -456
rect 257 -458 277 -456
rect 622 -456 642 -454
rect 576 -462 596 -460
rect 719 -460 721 -440
rect 729 -460 731 -440
rect 797 -457 799 -437
rect 827 -457 829 -437
rect 576 -472 596 -470
rect -33 -483 -13 -481
rect 330 -496 332 -476
rect 349 -496 351 -476
rect -102 -504 -82 -502
rect 122 -507 162 -505
rect 187 -507 227 -505
rect 409 -501 411 -481
rect 642 -487 662 -485
rect 446 -498 466 -496
rect 122 -517 162 -515
rect 187 -517 227 -515
rect -102 -534 -82 -532
rect 847 -477 849 -437
rect 857 -477 859 -437
rect 873 -477 875 -437
rect 883 -477 885 -437
rect 796 -483 816 -481
rect 557 -505 597 -503
rect 622 -505 662 -503
rect 865 -504 885 -502
rect 446 -508 466 -506
rect 557 -515 597 -513
rect 622 -515 662 -513
rect 122 -535 142 -533
rect -33 -555 -13 -553
rect -102 -599 -100 -559
rect -92 -599 -90 -559
rect -76 -599 -74 -559
rect -66 -599 -64 -559
rect 865 -534 885 -532
rect 188 -550 208 -548
rect -46 -599 -44 -579
rect -16 -599 -14 -579
rect 53 -580 55 -560
rect 63 -580 65 -560
rect 188 -560 208 -558
rect 142 -566 162 -564
rect 142 -576 162 -574
rect 188 -576 208 -574
rect 500 -579 502 -559
rect 519 -579 521 -559
rect 719 -580 721 -540
rect 729 -580 731 -540
rect 796 -555 816 -553
rect 633 -588 653 -586
rect 122 -607 162 -605
rect 211 -615 231 -613
rect 266 -615 286 -613
rect 122 -617 162 -615
rect 321 -620 341 -618
rect 122 -635 142 -633
rect 211 -634 231 -632
rect 409 -634 411 -594
rect 419 -634 421 -594
rect 797 -599 799 -579
rect 827 -599 829 -579
rect 847 -599 849 -559
rect 857 -599 859 -559
rect 873 -599 875 -559
rect 883 -599 885 -559
rect 452 -633 454 -613
rect 462 -633 464 -613
rect 478 -633 480 -613
rect 702 -609 722 -607
rect 519 -634 521 -614
rect 266 -639 286 -637
rect 321 -639 341 -637
rect 576 -646 578 -626
rect 633 -653 635 -613
rect 643 -653 645 -613
rect 659 -653 661 -613
rect 669 -653 671 -613
rect 689 -653 691 -633
rect 719 -653 721 -633
rect 763 -653 765 -633
rect 409 -699 411 -659
rect 419 -699 421 -659
rect 468 -679 470 -659
rect 478 -679 480 -659
rect 437 -699 439 -679
rect 509 -699 511 -659
rect 519 -699 521 -659
rect 537 -699 539 -679
rect 188 -745 190 -725
rect 232 -745 234 -725
rect 262 -745 264 -725
rect 282 -765 284 -725
rect 292 -765 294 -725
rect 308 -765 310 -725
rect 318 -765 320 -725
rect 576 -701 578 -681
rect 595 -701 597 -681
rect 343 -758 383 -756
rect 463 -758 483 -756
rect 343 -768 383 -766
rect 463 -768 483 -766
rect 231 -771 251 -769
rect 300 -792 320 -790
rect 356 -835 376 -833
rect 400 -852 402 -832
rect 472 -852 474 -832
rect 498 -835 518 -833
rect 356 -865 376 -863
rect 498 -865 518 -863
rect 356 -885 396 -883
rect 478 -885 518 -883
rect 356 -895 396 -893
rect 478 -895 518 -893
rect 356 -911 396 -909
rect 356 -921 396 -919
rect 421 -921 423 -901
rect 451 -921 453 -901
rect 478 -911 518 -909
rect 478 -921 518 -919
<< ndiffusion >>
rect 297 -92 303 -88
rect 293 -93 303 -92
rect 508 -92 514 -88
rect 508 -93 518 -92
rect 293 -97 303 -95
rect 293 -101 299 -97
rect 508 -97 518 -95
rect 512 -101 518 -97
rect 297 -118 303 -114
rect 293 -119 303 -118
rect 293 -123 303 -121
rect 293 -127 299 -123
rect 508 -118 514 -114
rect 508 -119 518 -118
rect 384 -131 389 -125
rect 388 -135 389 -131
rect 391 -129 392 -125
rect 391 -135 396 -129
rect 419 -129 420 -125
rect 415 -135 420 -129
rect 422 -131 427 -125
rect 508 -123 518 -121
rect 512 -127 518 -123
rect 422 -135 423 -131
rect 296 -148 312 -144
rect 292 -149 312 -148
rect 499 -148 515 -144
rect 499 -149 519 -148
rect 292 -153 312 -151
rect 296 -157 312 -153
rect 499 -153 519 -151
rect 292 -159 312 -157
rect 499 -157 515 -153
rect 292 -162 312 -161
rect 499 -159 519 -157
rect 499 -162 519 -161
rect 292 -166 308 -162
rect 296 -178 312 -174
rect 292 -179 312 -178
rect 292 -183 312 -181
rect 296 -187 312 -183
rect 503 -166 519 -162
rect 499 -178 515 -174
rect 499 -179 519 -178
rect 292 -189 312 -187
rect 292 -192 312 -191
rect 292 -196 308 -192
rect 499 -183 519 -181
rect 499 -187 515 -183
rect 499 -189 519 -187
rect 499 -192 519 -191
rect 363 -200 368 -194
rect 367 -204 368 -200
rect 370 -198 371 -194
rect 370 -204 375 -198
rect 440 -198 441 -194
rect 436 -204 441 -198
rect 443 -200 448 -194
rect 503 -196 519 -192
rect 443 -204 444 -200
rect 242 -221 248 -217
rect 242 -222 252 -221
rect 242 -225 252 -224
rect 246 -229 252 -225
rect 579 -237 580 -233
rect 173 -242 179 -238
rect 173 -243 183 -242
rect 575 -243 580 -237
rect 582 -239 588 -233
rect 582 -243 584 -239
rect 173 -246 183 -245
rect 177 -250 183 -246
rect 383 -251 399 -247
rect 383 -252 403 -251
rect 418 -251 424 -247
rect 414 -252 424 -251
rect 383 -262 403 -254
rect 414 -256 424 -254
rect 414 -260 420 -256
rect 414 -262 424 -260
rect 605 -237 606 -233
rect 601 -243 606 -237
rect 608 -239 614 -233
rect 608 -243 610 -239
rect 635 -236 636 -232
rect 631 -252 636 -236
rect 638 -236 640 -232
rect 644 -236 646 -232
rect 638 -252 646 -236
rect 648 -248 653 -232
rect 648 -252 649 -248
rect 665 -236 666 -232
rect 661 -252 666 -236
rect 668 -236 670 -232
rect 674 -236 676 -232
rect 668 -252 676 -236
rect 678 -248 683 -232
rect 678 -252 679 -248
rect 709 -246 710 -242
rect 705 -252 710 -246
rect 712 -248 717 -242
rect 712 -252 713 -248
rect 383 -265 403 -264
rect 387 -269 403 -265
rect 414 -265 424 -264
rect 418 -269 424 -265
rect 151 -305 152 -301
rect 73 -312 79 -308
rect 147 -311 152 -305
rect 154 -307 159 -301
rect 154 -311 155 -307
rect 185 -305 186 -301
rect 69 -313 79 -312
rect 69 -316 79 -315
rect 69 -320 75 -316
rect 181 -321 186 -305
rect 188 -317 196 -301
rect 188 -321 190 -317
rect 194 -321 196 -317
rect 198 -317 203 -301
rect 198 -321 199 -317
rect 215 -305 216 -301
rect 211 -321 216 -305
rect 218 -317 226 -301
rect 218 -321 220 -317
rect 224 -321 226 -317
rect 228 -317 233 -301
rect 228 -321 229 -317
rect 142 -333 148 -329
rect 138 -334 148 -333
rect 138 -337 148 -336
rect 138 -341 144 -337
rect 254 -314 256 -310
rect 250 -320 256 -314
rect 258 -316 263 -310
rect 258 -320 259 -316
rect 280 -314 282 -310
rect 276 -320 282 -314
rect 284 -316 289 -310
rect 284 -320 285 -316
rect 790 -265 796 -261
rect 786 -266 796 -265
rect 786 -269 796 -268
rect 786 -273 792 -269
rect 859 -286 865 -282
rect 855 -287 865 -286
rect 681 -307 687 -303
rect 681 -308 691 -307
rect 681 -311 691 -310
rect 685 -315 691 -311
rect 612 -328 618 -324
rect 612 -329 622 -328
rect 341 -336 342 -332
rect 337 -352 342 -336
rect 344 -352 352 -332
rect 354 -348 359 -332
rect 354 -352 355 -348
rect 382 -347 383 -343
rect 378 -353 383 -347
rect 385 -349 390 -343
rect 385 -353 386 -349
rect 396 -356 401 -350
rect 400 -360 401 -356
rect 403 -354 405 -350
rect 409 -354 411 -350
rect 403 -360 411 -354
rect 413 -356 418 -350
rect 612 -332 622 -331
rect 616 -336 622 -332
rect 855 -290 865 -289
rect 855 -294 861 -290
rect 413 -360 414 -356
rect 666 -358 682 -354
rect 662 -359 682 -358
rect 749 -360 754 -354
rect 293 -371 299 -367
rect 289 -372 299 -371
rect 475 -370 476 -366
rect 289 -375 299 -374
rect 293 -379 299 -375
rect 471 -376 476 -370
rect 478 -372 483 -366
rect 662 -369 682 -361
rect 753 -364 754 -360
rect 756 -358 758 -354
rect 756 -364 762 -358
rect 478 -376 479 -372
rect 662 -372 682 -371
rect 662 -376 678 -372
rect -103 -410 -102 -406
rect -107 -416 -102 -410
rect -100 -412 -94 -406
rect -100 -416 -98 -412
rect -77 -410 -76 -406
rect -81 -416 -76 -410
rect -74 -412 -68 -406
rect -74 -416 -72 -412
rect -47 -409 -46 -405
rect -51 -425 -46 -409
rect -44 -409 -42 -405
rect -38 -409 -36 -405
rect -44 -425 -36 -409
rect -34 -421 -29 -405
rect -34 -425 -33 -421
rect -17 -409 -16 -405
rect -21 -425 -16 -409
rect -14 -409 -12 -405
rect -8 -409 -6 -405
rect -14 -425 -6 -409
rect -4 -421 1 -405
rect 32 -407 37 -401
rect 36 -411 37 -407
rect 39 -405 41 -401
rect 39 -411 45 -405
rect -4 -425 -3 -421
rect 58 -407 63 -401
rect 62 -411 63 -407
rect 65 -405 67 -401
rect 65 -411 71 -405
rect 239 -390 245 -386
rect 235 -391 245 -390
rect 293 -390 299 -386
rect 534 -380 540 -376
rect 534 -381 544 -380
rect 775 -360 780 -354
rect 779 -364 780 -360
rect 782 -358 784 -354
rect 782 -364 788 -358
rect 805 -361 810 -345
rect 809 -365 810 -361
rect 812 -361 820 -345
rect 812 -365 814 -361
rect 818 -365 820 -361
rect 822 -349 823 -345
rect 822 -365 827 -349
rect 835 -361 840 -345
rect 839 -365 840 -361
rect 842 -361 850 -345
rect 842 -365 844 -361
rect 848 -365 850 -361
rect 852 -349 853 -345
rect 852 -365 857 -349
rect 879 -351 884 -345
rect 883 -355 884 -351
rect 886 -349 887 -345
rect 886 -355 891 -349
rect 534 -384 544 -383
rect 538 -388 544 -384
rect 289 -391 299 -390
rect 88 -408 93 -392
rect 92 -412 93 -408
rect 95 -408 103 -392
rect 95 -412 97 -408
rect 101 -412 103 -408
rect 105 -396 106 -392
rect 105 -412 110 -396
rect 118 -408 123 -392
rect 122 -412 123 -408
rect 125 -408 133 -392
rect 125 -412 127 -408
rect 131 -412 133 -408
rect 135 -396 136 -392
rect 135 -412 140 -396
rect 235 -394 245 -393
rect 235 -398 241 -394
rect 289 -394 299 -393
rect 289 -398 295 -394
rect 531 -398 537 -394
rect 527 -399 537 -398
rect 527 -403 537 -401
rect 527 -407 533 -403
rect 527 -409 537 -407
rect 681 -402 687 -398
rect 681 -403 691 -402
rect 527 -412 537 -411
rect 531 -416 537 -412
rect 681 -407 691 -405
rect 685 -411 691 -407
rect 681 -413 691 -411
rect 681 -416 691 -415
rect 681 -420 687 -416
rect 293 -436 299 -432
rect 289 -437 299 -436
rect -1 -480 5 -476
rect 289 -440 299 -439
rect 293 -444 299 -440
rect 456 -424 457 -420
rect 452 -430 457 -424
rect 459 -424 460 -420
rect 459 -430 464 -424
rect 475 -424 476 -420
rect 471 -430 476 -424
rect 478 -426 483 -420
rect 782 -421 787 -405
rect 786 -425 787 -421
rect 789 -409 791 -405
rect 795 -409 797 -405
rect 789 -425 797 -409
rect 799 -409 800 -405
rect 799 -425 804 -409
rect 812 -421 817 -405
rect 816 -425 817 -421
rect 819 -409 821 -405
rect 825 -409 827 -405
rect 819 -425 827 -409
rect 829 -409 830 -405
rect 829 -425 834 -409
rect 478 -430 479 -426
rect 239 -455 245 -451
rect 235 -456 245 -455
rect 293 -455 299 -451
rect 554 -443 560 -439
rect 554 -444 564 -443
rect 666 -443 682 -439
rect 851 -412 857 -406
rect 855 -416 857 -412
rect 859 -410 860 -406
rect 859 -416 864 -410
rect 877 -412 883 -406
rect 881 -416 883 -412
rect 885 -410 886 -406
rect 885 -416 890 -410
rect 662 -444 682 -443
rect 554 -447 564 -446
rect 558 -451 564 -447
rect 662 -454 682 -446
rect 289 -456 299 -455
rect 348 -458 349 -454
rect 235 -459 245 -458
rect 235 -463 241 -459
rect 289 -459 299 -458
rect 289 -463 295 -459
rect 344 -464 349 -458
rect 351 -460 356 -454
rect 536 -459 552 -455
rect 536 -460 556 -459
rect 351 -464 352 -460
rect 662 -457 682 -456
rect 662 -461 678 -457
rect 536 -470 556 -462
rect 536 -473 556 -472
rect -1 -481 9 -480
rect -1 -484 9 -483
rect 3 -488 9 -484
rect -70 -501 -64 -497
rect 540 -477 556 -473
rect 778 -480 784 -476
rect -70 -502 -60 -501
rect -70 -505 -60 -504
rect -66 -509 -60 -505
rect 48 -505 53 -499
rect 52 -509 53 -505
rect 55 -503 57 -499
rect 61 -503 63 -499
rect 55 -509 63 -503
rect 65 -505 70 -499
rect 97 -504 103 -500
rect 93 -505 103 -504
rect 246 -504 252 -500
rect 246 -505 256 -504
rect 65 -509 66 -505
rect 93 -509 103 -507
rect 93 -513 99 -509
rect 93 -515 103 -513
rect 246 -509 256 -507
rect 678 -484 684 -480
rect 674 -485 684 -484
rect 718 -484 719 -480
rect 490 -495 506 -491
rect 674 -488 684 -487
rect 674 -492 680 -488
rect 486 -496 506 -495
rect 250 -513 256 -509
rect 246 -515 256 -513
rect 329 -512 330 -508
rect 93 -518 103 -517
rect 52 -524 53 -520
rect -66 -531 -60 -527
rect -70 -532 -60 -531
rect -70 -535 -60 -534
rect -70 -539 -64 -535
rect 48 -540 53 -524
rect 55 -540 63 -520
rect 65 -536 70 -520
rect 97 -522 103 -518
rect 246 -518 256 -517
rect 325 -518 330 -512
rect 332 -512 333 -508
rect 332 -518 337 -512
rect 348 -512 349 -508
rect 344 -518 349 -512
rect 351 -514 356 -508
rect 486 -506 506 -498
rect 532 -502 538 -498
rect 528 -503 538 -502
rect 681 -502 687 -498
rect 714 -500 719 -484
rect 721 -500 729 -480
rect 731 -496 736 -480
rect 774 -481 784 -480
rect 774 -484 784 -483
rect 774 -488 780 -484
rect 731 -500 732 -496
rect 681 -503 691 -502
rect 847 -501 853 -497
rect 843 -502 853 -501
rect 843 -505 853 -504
rect 528 -507 538 -505
rect 486 -509 506 -508
rect 486 -513 502 -509
rect 528 -511 534 -507
rect 528 -513 538 -511
rect 681 -507 691 -505
rect 685 -511 691 -507
rect 843 -509 849 -505
rect 681 -513 691 -511
rect 351 -518 352 -514
rect 246 -522 252 -518
rect 404 -519 409 -513
rect 408 -523 409 -519
rect 411 -517 412 -513
rect 718 -515 719 -511
rect 411 -523 416 -517
rect 528 -516 538 -515
rect 532 -520 538 -516
rect 681 -516 691 -515
rect 681 -520 687 -516
rect 714 -521 719 -515
rect 721 -517 729 -511
rect 721 -521 723 -517
rect 727 -521 729 -517
rect 731 -515 732 -511
rect 731 -521 736 -515
rect 104 -532 110 -528
rect 100 -533 110 -532
rect 65 -540 66 -536
rect 100 -536 110 -535
rect 100 -540 106 -536
rect 3 -552 9 -548
rect -1 -553 9 -552
rect -1 -556 9 -555
rect -1 -560 5 -556
rect 495 -543 500 -537
rect 228 -547 244 -543
rect 499 -547 500 -543
rect 502 -543 507 -537
rect 502 -547 503 -543
rect 514 -543 519 -537
rect 518 -547 519 -543
rect 521 -541 522 -537
rect 843 -531 849 -527
rect 843 -532 853 -531
rect 843 -535 853 -534
rect 847 -539 853 -535
rect 521 -547 526 -541
rect 228 -548 248 -547
rect 228 -558 248 -550
rect 106 -563 122 -559
rect 102 -564 122 -563
rect 228 -561 248 -560
rect 232 -565 248 -561
rect 102 -574 122 -566
rect 408 -569 409 -565
rect 220 -573 226 -569
rect 220 -574 230 -573
rect 404 -575 409 -569
rect 411 -571 419 -565
rect 411 -575 413 -571
rect 417 -575 419 -571
rect 421 -569 422 -565
rect 421 -575 426 -569
rect 102 -577 122 -576
rect 102 -581 118 -577
rect 220 -577 230 -576
rect 224 -581 230 -577
rect 451 -577 452 -573
rect 447 -593 452 -577
rect 454 -593 462 -573
rect 464 -589 469 -573
rect 464 -593 465 -589
rect 774 -552 780 -548
rect 774 -553 784 -552
rect 774 -556 784 -555
rect 778 -560 784 -556
rect 669 -585 675 -581
rect 665 -586 675 -585
rect -107 -626 -102 -620
rect -103 -630 -102 -626
rect -100 -624 -98 -620
rect -100 -630 -94 -624
rect -81 -626 -76 -620
rect -77 -630 -76 -626
rect -74 -624 -72 -620
rect -74 -630 -68 -624
rect 97 -604 103 -600
rect 93 -605 103 -604
rect 93 -609 103 -607
rect -51 -627 -46 -611
rect -47 -631 -46 -627
rect -44 -627 -36 -611
rect -44 -631 -42 -627
rect -38 -631 -36 -627
rect -34 -615 -33 -611
rect -34 -631 -29 -615
rect -21 -627 -16 -611
rect -17 -631 -16 -627
rect -14 -627 -6 -611
rect -14 -631 -12 -627
rect -8 -631 -6 -627
rect -4 -615 -3 -611
rect 93 -613 99 -609
rect 93 -615 103 -613
rect 193 -612 199 -608
rect 189 -613 199 -612
rect 247 -612 253 -608
rect 243 -613 253 -612
rect -4 -631 1 -615
rect 189 -616 199 -615
rect 93 -618 103 -617
rect 97 -622 103 -618
rect 189 -620 195 -616
rect 243 -616 253 -615
rect 243 -620 249 -616
rect 357 -617 363 -613
rect 353 -618 363 -617
rect 353 -621 363 -620
rect 357 -625 363 -621
rect 104 -632 110 -628
rect 100 -633 110 -632
rect 189 -631 195 -627
rect 189 -632 199 -631
rect 100 -636 110 -635
rect 100 -640 106 -636
rect 189 -635 199 -634
rect 189 -639 195 -635
rect 303 -636 309 -632
rect 299 -637 309 -636
rect 357 -636 363 -632
rect 477 -595 478 -591
rect 473 -601 478 -595
rect 480 -597 485 -591
rect 480 -601 481 -597
rect 514 -597 519 -591
rect 518 -601 519 -597
rect 521 -595 522 -591
rect 665 -589 675 -588
rect 665 -593 671 -589
rect 521 -601 526 -595
rect 738 -606 744 -602
rect 734 -607 744 -606
rect 353 -637 363 -636
rect 299 -640 309 -639
rect 299 -644 305 -640
rect 353 -640 363 -639
rect 353 -644 359 -640
rect 734 -610 744 -609
rect 734 -614 740 -610
rect 786 -615 787 -611
rect 782 -631 787 -615
rect 789 -627 797 -611
rect 789 -631 791 -627
rect 795 -631 797 -627
rect 799 -627 804 -611
rect 799 -631 800 -627
rect 816 -615 817 -611
rect 812 -631 817 -615
rect 819 -627 827 -611
rect 819 -631 821 -627
rect 825 -631 827 -627
rect 829 -627 834 -611
rect 829 -631 830 -627
rect 855 -624 857 -620
rect 851 -630 857 -624
rect 859 -626 864 -620
rect 859 -630 860 -626
rect 881 -624 883 -620
rect 877 -630 883 -624
rect 885 -626 890 -620
rect 885 -630 886 -626
rect 183 -709 188 -703
rect 187 -713 188 -709
rect 190 -707 191 -703
rect 190 -713 195 -707
rect 217 -709 222 -693
rect 221 -713 222 -709
rect 224 -697 226 -693
rect 230 -697 232 -693
rect 224 -713 232 -697
rect 234 -697 235 -693
rect 234 -713 239 -697
rect 247 -709 252 -693
rect 251 -713 252 -709
rect 254 -697 256 -693
rect 260 -697 262 -693
rect 254 -713 262 -697
rect 264 -697 265 -693
rect 264 -713 269 -697
rect 286 -700 292 -694
rect 290 -704 292 -700
rect 294 -698 295 -694
rect 294 -704 299 -698
rect 312 -700 318 -694
rect 316 -704 318 -700
rect 320 -698 321 -694
rect 320 -704 325 -698
rect 571 -665 576 -659
rect 575 -669 576 -665
rect 578 -663 579 -659
rect 578 -669 583 -663
rect 628 -680 633 -674
rect 432 -717 437 -711
rect 404 -724 409 -718
rect 213 -768 219 -764
rect 209 -769 219 -768
rect 408 -728 409 -724
rect 411 -722 413 -718
rect 417 -722 419 -718
rect 411 -728 419 -722
rect 421 -724 426 -718
rect 436 -721 437 -717
rect 439 -715 440 -711
rect 439 -721 444 -715
rect 463 -715 468 -699
rect 467 -719 468 -715
rect 470 -719 478 -699
rect 480 -703 481 -699
rect 480 -719 485 -703
rect 632 -684 633 -680
rect 635 -678 637 -674
rect 635 -684 641 -678
rect 532 -717 537 -711
rect 421 -728 422 -724
rect 504 -724 509 -718
rect 508 -728 509 -724
rect 511 -722 513 -718
rect 517 -722 519 -718
rect 511 -728 519 -722
rect 521 -724 526 -718
rect 536 -721 537 -717
rect 539 -715 540 -711
rect 654 -680 659 -674
rect 658 -684 659 -680
rect 661 -678 663 -674
rect 661 -684 667 -678
rect 684 -681 689 -665
rect 688 -685 689 -681
rect 691 -681 699 -665
rect 691 -685 693 -681
rect 697 -685 699 -681
rect 701 -669 702 -665
rect 701 -685 706 -669
rect 714 -681 719 -665
rect 718 -685 719 -681
rect 721 -681 729 -665
rect 721 -685 723 -681
rect 727 -685 729 -681
rect 731 -669 732 -665
rect 731 -685 736 -669
rect 758 -671 763 -665
rect 762 -675 763 -671
rect 765 -669 766 -665
rect 765 -675 770 -669
rect 539 -721 544 -715
rect 571 -719 576 -713
rect 521 -728 522 -724
rect 575 -723 576 -719
rect 578 -717 579 -713
rect 578 -723 583 -717
rect 594 -717 595 -713
rect 590 -723 595 -717
rect 597 -717 598 -713
rect 597 -723 602 -717
rect 402 -755 408 -751
rect 402 -756 412 -755
rect 423 -755 439 -751
rect 423 -756 443 -755
rect 402 -760 412 -758
rect 406 -764 412 -760
rect 402 -766 412 -764
rect 423 -766 443 -758
rect 209 -772 219 -771
rect 209 -776 215 -772
rect 402 -769 412 -768
rect 402 -773 408 -769
rect 423 -769 443 -768
rect 427 -773 443 -769
rect 282 -789 288 -785
rect 278 -790 288 -789
rect 278 -793 288 -792
rect 278 -797 284 -793
rect 399 -814 400 -810
rect 324 -822 340 -818
rect 395 -820 400 -814
rect 402 -816 407 -810
rect 402 -820 403 -816
rect 467 -816 472 -810
rect 471 -820 472 -816
rect 474 -814 475 -810
rect 474 -820 479 -814
rect 324 -823 344 -822
rect 324 -827 344 -825
rect 328 -831 344 -827
rect 324 -833 344 -831
rect 534 -822 550 -818
rect 530 -823 550 -822
rect 530 -827 550 -825
rect 324 -836 344 -835
rect 328 -840 344 -836
rect 324 -852 340 -848
rect 530 -831 546 -827
rect 530 -833 550 -831
rect 530 -836 550 -835
rect 530 -840 546 -836
rect 534 -852 550 -848
rect 324 -853 344 -852
rect 324 -857 344 -855
rect 530 -853 550 -852
rect 328 -861 344 -857
rect 530 -857 550 -855
rect 324 -863 344 -861
rect 530 -861 546 -857
rect 530 -863 550 -861
rect 324 -866 344 -865
rect 328 -870 344 -866
rect 530 -866 550 -865
rect 530 -870 546 -866
rect 420 -883 421 -879
rect 325 -891 331 -887
rect 325 -893 335 -891
rect 416 -889 421 -883
rect 423 -885 428 -879
rect 423 -889 424 -885
rect 446 -885 451 -879
rect 450 -889 451 -885
rect 453 -883 454 -879
rect 453 -889 458 -883
rect 325 -896 335 -895
rect 329 -900 335 -896
rect 543 -891 549 -887
rect 539 -893 549 -891
rect 539 -896 549 -895
rect 539 -900 545 -896
rect 325 -917 331 -913
rect 325 -919 335 -917
rect 543 -917 549 -913
rect 539 -919 549 -917
rect 325 -922 335 -921
rect 329 -926 335 -922
rect 539 -922 549 -921
rect 539 -926 545 -922
<< pdiffusion >>
rect 324 -92 360 -88
rect 324 -93 364 -92
rect 451 -92 487 -88
rect 447 -93 487 -92
rect 324 -97 364 -95
rect 328 -101 364 -97
rect 324 -103 364 -101
rect 388 -97 389 -93
rect 324 -106 364 -105
rect 328 -110 364 -106
rect 384 -113 389 -97
rect 391 -109 396 -93
rect 391 -113 392 -109
rect 415 -109 420 -93
rect 419 -113 420 -109
rect 422 -97 423 -93
rect 422 -113 427 -97
rect 447 -97 487 -95
rect 447 -101 483 -97
rect 447 -103 487 -101
rect 447 -106 487 -105
rect 447 -110 483 -106
rect 324 -118 360 -114
rect 324 -119 364 -118
rect 324 -123 364 -121
rect 324 -127 360 -123
rect 451 -118 487 -114
rect 447 -119 487 -118
rect 447 -123 487 -121
rect 324 -129 364 -127
rect 324 -132 364 -131
rect 328 -136 360 -132
rect 451 -127 487 -123
rect 447 -129 487 -127
rect 447 -132 487 -131
rect 451 -136 483 -132
rect 324 -148 340 -144
rect 324 -149 344 -148
rect 471 -148 487 -144
rect 467 -149 487 -148
rect 324 -152 344 -151
rect 328 -156 344 -152
rect 467 -152 487 -151
rect 467 -156 483 -152
rect 367 -166 368 -162
rect 324 -178 340 -174
rect 324 -179 344 -178
rect 324 -182 344 -181
rect 363 -182 368 -166
rect 370 -178 375 -162
rect 370 -182 371 -178
rect 436 -178 441 -162
rect 440 -182 441 -178
rect 443 -166 444 -162
rect 443 -182 448 -166
rect 471 -178 487 -174
rect 467 -179 487 -178
rect 467 -182 487 -181
rect 328 -186 344 -182
rect 467 -186 483 -182
rect 268 -221 284 -217
rect 264 -222 284 -221
rect 264 -225 284 -224
rect 264 -229 280 -225
rect 199 -242 215 -238
rect 195 -243 215 -242
rect 195 -246 215 -245
rect 195 -250 211 -246
rect 245 -253 246 -249
rect 147 -285 152 -269
rect 151 -289 152 -285
rect 154 -273 155 -269
rect 154 -289 159 -273
rect 191 -285 196 -269
rect 195 -289 196 -285
rect 198 -273 199 -269
rect 198 -289 203 -273
rect 221 -285 226 -269
rect 225 -289 226 -285
rect 228 -273 229 -269
rect 228 -289 233 -273
rect 241 -285 246 -253
rect 245 -289 246 -285
rect 248 -253 250 -249
rect 254 -253 256 -249
rect 248 -289 256 -253
rect 258 -253 259 -249
rect 258 -289 263 -253
rect 267 -285 272 -249
rect 271 -289 272 -285
rect 274 -285 282 -249
rect 274 -289 276 -285
rect 280 -289 282 -285
rect 284 -253 285 -249
rect 347 -251 363 -247
rect 343 -252 363 -251
rect 443 -251 479 -247
rect 443 -252 483 -251
rect 284 -289 289 -253
rect 343 -256 363 -254
rect 343 -260 359 -256
rect 343 -262 363 -260
rect 443 -262 483 -254
rect 343 -265 363 -264
rect 347 -269 363 -265
rect 443 -265 483 -264
rect 447 -269 483 -265
rect 37 -312 53 -308
rect 37 -313 57 -312
rect 37 -316 57 -315
rect 41 -320 57 -316
rect 106 -333 122 -329
rect 106 -334 126 -333
rect 106 -337 126 -336
rect 36 -344 37 -340
rect 32 -380 37 -344
rect 39 -376 47 -340
rect 39 -380 41 -376
rect 45 -380 47 -376
rect 49 -376 54 -340
rect 49 -380 50 -376
rect 62 -344 63 -340
rect 58 -380 63 -344
rect 65 -344 67 -340
rect 71 -344 73 -340
rect 65 -380 73 -344
rect 75 -344 76 -340
rect 110 -341 126 -337
rect 341 -296 342 -292
rect 337 -312 342 -296
rect 344 -308 352 -292
rect 344 -312 346 -308
rect 350 -312 352 -308
rect 354 -296 355 -292
rect 354 -312 359 -296
rect 378 -327 383 -311
rect 382 -331 383 -327
rect 385 -315 386 -311
rect 385 -331 390 -315
rect 396 -327 401 -291
rect 400 -331 401 -327
rect 403 -331 411 -291
rect 413 -295 414 -291
rect 413 -331 418 -295
rect 575 -300 580 -264
rect 579 -304 580 -300
rect 582 -268 584 -264
rect 588 -268 590 -264
rect 582 -304 590 -268
rect 592 -268 593 -264
rect 592 -304 597 -268
rect 601 -300 606 -264
rect 605 -304 606 -300
rect 608 -300 616 -264
rect 608 -304 610 -300
rect 614 -304 616 -300
rect 618 -268 619 -264
rect 618 -300 623 -268
rect 631 -280 636 -264
rect 635 -284 636 -280
rect 638 -268 639 -264
rect 638 -284 643 -268
rect 661 -280 666 -264
rect 665 -284 666 -280
rect 668 -268 669 -264
rect 668 -284 673 -268
rect 705 -280 710 -264
rect 709 -284 710 -280
rect 712 -268 713 -264
rect 754 -265 770 -261
rect 754 -266 774 -265
rect 712 -284 717 -268
rect 754 -269 774 -268
rect 758 -273 774 -269
rect 823 -286 839 -282
rect 823 -287 843 -286
rect 823 -290 843 -289
rect 618 -304 619 -300
rect 753 -297 754 -293
rect 653 -307 669 -303
rect 649 -308 669 -307
rect 649 -311 669 -310
rect 649 -315 665 -311
rect 584 -328 600 -324
rect 580 -329 600 -328
rect 75 -376 80 -344
rect 580 -332 600 -331
rect 471 -349 476 -333
rect 475 -353 476 -349
rect 478 -337 479 -333
rect 580 -336 596 -332
rect 749 -333 754 -297
rect 756 -329 764 -293
rect 756 -333 758 -329
rect 762 -333 764 -329
rect 766 -329 771 -293
rect 766 -333 767 -329
rect 779 -297 780 -293
rect 775 -333 780 -297
rect 782 -297 784 -293
rect 788 -297 790 -293
rect 782 -333 790 -297
rect 792 -297 793 -293
rect 827 -294 843 -290
rect 792 -329 797 -297
rect 792 -333 793 -329
rect 809 -317 810 -313
rect 805 -333 810 -317
rect 812 -329 817 -313
rect 812 -333 813 -329
rect 839 -317 840 -313
rect 835 -333 840 -317
rect 842 -329 847 -313
rect 842 -333 843 -329
rect 883 -317 884 -313
rect 879 -333 884 -317
rect 886 -329 891 -313
rect 886 -333 887 -329
rect 478 -353 483 -337
rect 75 -380 76 -376
rect 92 -364 93 -360
rect 88 -380 93 -364
rect 95 -376 100 -360
rect 95 -380 96 -376
rect 122 -364 123 -360
rect 118 -380 123 -364
rect 125 -376 130 -360
rect 626 -358 642 -354
rect 622 -359 642 -358
rect 622 -363 642 -361
rect 257 -371 273 -367
rect 257 -372 277 -371
rect 125 -380 126 -376
rect 257 -375 277 -374
rect 257 -379 273 -375
rect 622 -367 638 -363
rect 622 -369 642 -367
rect 622 -372 642 -371
rect 626 -376 642 -372
rect 202 -390 218 -386
rect 202 -391 222 -390
rect 257 -390 273 -386
rect 257 -391 277 -390
rect 560 -380 576 -376
rect 556 -381 576 -380
rect 556 -384 576 -383
rect 556 -388 572 -384
rect 202 -394 222 -393
rect 206 -398 222 -394
rect 257 -394 277 -393
rect 261 -398 277 -394
rect 452 -404 457 -388
rect 456 -408 457 -404
rect 459 -404 464 -388
rect 459 -408 460 -404
rect 471 -404 476 -388
rect 475 -408 476 -404
rect 478 -392 479 -388
rect 478 -408 483 -392
rect 560 -398 596 -394
rect 556 -399 596 -398
rect 556 -409 596 -401
rect 622 -402 658 -398
rect 622 -403 662 -402
rect 556 -412 596 -411
rect 556 -416 592 -412
rect 622 -413 662 -405
rect 622 -416 662 -415
rect 626 -420 662 -416
rect 257 -436 273 -432
rect 257 -437 277 -436
rect 344 -437 349 -421
rect -107 -473 -102 -437
rect -103 -477 -102 -473
rect -100 -441 -98 -437
rect -94 -441 -92 -437
rect -100 -477 -92 -441
rect -90 -441 -89 -437
rect -90 -477 -85 -441
rect -81 -473 -76 -437
rect -77 -477 -76 -473
rect -74 -473 -66 -437
rect -74 -477 -72 -473
rect -68 -477 -66 -473
rect -64 -441 -63 -437
rect -64 -473 -59 -441
rect -51 -453 -46 -437
rect -47 -457 -46 -453
rect -44 -441 -43 -437
rect -44 -457 -39 -441
rect -21 -453 -16 -437
rect -17 -457 -16 -453
rect -14 -441 -13 -437
rect -14 -457 -9 -441
rect -64 -477 -63 -473
rect 48 -476 53 -440
rect -29 -480 -13 -476
rect -33 -481 -13 -480
rect 52 -480 53 -476
rect 55 -480 63 -440
rect 65 -476 70 -440
rect 257 -440 277 -439
rect 257 -444 273 -440
rect 348 -441 349 -437
rect 351 -425 352 -421
rect 351 -441 356 -425
rect 202 -455 218 -451
rect 202 -456 222 -455
rect 257 -455 273 -451
rect 257 -456 277 -455
rect 580 -443 596 -439
rect 576 -444 596 -443
rect 626 -443 642 -439
rect 622 -444 642 -443
rect 718 -444 719 -440
rect 576 -447 596 -446
rect 576 -451 592 -447
rect 622 -448 642 -446
rect 622 -452 638 -448
rect 622 -454 642 -452
rect 202 -459 222 -458
rect 206 -463 222 -459
rect 257 -459 277 -458
rect 261 -463 277 -459
rect 576 -459 592 -455
rect 576 -460 596 -459
rect 622 -457 642 -456
rect 626 -461 642 -457
rect 714 -460 719 -444
rect 721 -456 729 -440
rect 721 -460 723 -456
rect 727 -460 729 -456
rect 731 -444 732 -440
rect 731 -460 736 -444
rect 796 -441 797 -437
rect 792 -457 797 -441
rect 799 -453 804 -437
rect 799 -457 800 -453
rect 826 -441 827 -437
rect 822 -457 827 -441
rect 829 -453 834 -437
rect 829 -457 830 -453
rect 846 -441 847 -437
rect 576 -464 596 -462
rect 580 -468 596 -464
rect 576 -470 596 -468
rect 65 -480 66 -476
rect -33 -484 -13 -483
rect -33 -488 -17 -484
rect -98 -501 -82 -497
rect -102 -502 -82 -501
rect 325 -492 330 -476
rect 329 -496 330 -492
rect 332 -492 337 -476
rect 332 -496 333 -492
rect 344 -492 349 -476
rect 348 -496 349 -492
rect 351 -480 352 -476
rect 576 -473 596 -472
rect 576 -477 592 -473
rect 351 -496 356 -480
rect 842 -473 847 -441
rect 408 -485 409 -481
rect -102 -505 -82 -504
rect -102 -509 -86 -505
rect 122 -504 158 -500
rect 122 -505 162 -504
rect 191 -504 227 -500
rect 187 -505 227 -504
rect 122 -515 162 -507
rect 187 -515 227 -507
rect 404 -501 409 -485
rect 411 -497 416 -481
rect 642 -484 658 -480
rect 642 -485 662 -484
rect 642 -488 662 -487
rect 450 -495 466 -491
rect 446 -496 466 -495
rect 646 -492 662 -488
rect 411 -501 412 -497
rect 446 -500 466 -498
rect -102 -531 -86 -527
rect -102 -532 -82 -531
rect -102 -535 -82 -534
rect -98 -539 -82 -535
rect 122 -518 162 -517
rect 126 -522 162 -518
rect 187 -518 227 -517
rect 187 -522 223 -518
rect 446 -504 462 -500
rect 446 -506 466 -504
rect 561 -502 597 -498
rect 557 -503 597 -502
rect 622 -502 658 -498
rect 622 -503 662 -502
rect 796 -480 812 -476
rect 846 -477 847 -473
rect 849 -473 857 -437
rect 849 -477 851 -473
rect 855 -477 857 -473
rect 859 -473 864 -437
rect 859 -477 860 -473
rect 872 -441 873 -437
rect 868 -477 873 -441
rect 875 -441 877 -437
rect 881 -441 883 -437
rect 875 -477 883 -441
rect 885 -473 890 -437
rect 885 -477 886 -473
rect 796 -481 816 -480
rect 796 -484 816 -483
rect 800 -488 816 -484
rect 865 -501 881 -497
rect 865 -502 885 -501
rect 446 -509 466 -508
rect 450 -513 466 -509
rect 557 -513 597 -505
rect 622 -513 662 -505
rect 865 -505 885 -504
rect 869 -509 885 -505
rect 557 -516 597 -515
rect 557 -520 571 -516
rect 575 -520 593 -516
rect 622 -516 662 -515
rect 626 -520 662 -516
rect 122 -532 138 -528
rect 122 -533 142 -532
rect 122 -536 142 -535
rect 126 -540 142 -536
rect -33 -552 -17 -548
rect -33 -553 -13 -552
rect -33 -556 -13 -555
rect -103 -563 -102 -559
rect -107 -599 -102 -563
rect -100 -595 -92 -559
rect -100 -599 -98 -595
rect -94 -599 -92 -595
rect -90 -595 -85 -559
rect -90 -599 -89 -595
rect -77 -563 -76 -559
rect -81 -599 -76 -563
rect -74 -563 -72 -559
rect -68 -563 -66 -559
rect -74 -599 -66 -563
rect -64 -563 -63 -559
rect -29 -560 -13 -556
rect 192 -547 208 -543
rect 188 -548 208 -547
rect 869 -531 885 -527
rect 865 -532 885 -531
rect 865 -535 885 -534
rect 865 -539 881 -535
rect 718 -544 719 -540
rect 188 -552 208 -550
rect 188 -556 204 -552
rect 188 -558 208 -556
rect -64 -595 -59 -563
rect 48 -576 53 -560
rect -64 -599 -63 -595
rect -47 -583 -46 -579
rect -51 -599 -46 -583
rect -44 -595 -39 -579
rect -44 -599 -43 -595
rect -17 -583 -16 -579
rect -21 -599 -16 -583
rect -14 -595 -9 -579
rect 52 -580 53 -576
rect 55 -564 57 -560
rect 61 -564 63 -560
rect 55 -580 63 -564
rect 65 -576 70 -560
rect 142 -563 158 -559
rect 142 -564 162 -563
rect 188 -561 208 -560
rect 192 -565 208 -561
rect 499 -563 500 -559
rect 142 -568 162 -566
rect 146 -572 162 -568
rect 142 -574 162 -572
rect 192 -573 208 -569
rect 188 -574 208 -573
rect 65 -580 66 -576
rect 142 -577 162 -576
rect 142 -581 158 -577
rect 188 -577 208 -576
rect 188 -581 204 -577
rect 495 -579 500 -563
rect 502 -563 503 -559
rect 502 -579 507 -563
rect 518 -563 519 -559
rect 514 -579 519 -563
rect 521 -575 526 -559
rect 521 -579 522 -575
rect 714 -580 719 -544
rect 721 -580 729 -540
rect 731 -544 732 -540
rect 731 -580 736 -544
rect 800 -552 816 -548
rect 796 -553 816 -552
rect 796 -556 816 -555
rect 796 -560 812 -556
rect 846 -563 847 -559
rect 633 -585 649 -581
rect 633 -586 653 -585
rect 633 -589 653 -588
rect -14 -599 -13 -595
rect 122 -604 158 -600
rect 122 -605 162 -604
rect 122 -615 162 -607
rect 211 -612 227 -608
rect 211 -613 231 -612
rect 266 -612 282 -608
rect 266 -613 286 -612
rect 122 -618 162 -617
rect 126 -622 162 -618
rect 211 -616 231 -615
rect 215 -620 231 -616
rect 266 -616 286 -615
rect 270 -620 286 -616
rect 321 -617 337 -613
rect 321 -618 341 -617
rect 321 -621 341 -620
rect 321 -625 337 -621
rect 122 -632 138 -628
rect 215 -631 231 -627
rect 211 -632 231 -631
rect 404 -630 409 -594
rect 122 -633 142 -632
rect 122 -636 142 -635
rect 126 -640 142 -636
rect 211 -635 231 -634
rect 215 -639 231 -635
rect 266 -636 282 -632
rect 266 -637 286 -636
rect 321 -636 337 -632
rect 321 -637 341 -636
rect 408 -634 409 -630
rect 411 -634 419 -594
rect 421 -598 422 -594
rect 421 -634 426 -598
rect 637 -593 653 -589
rect 792 -595 797 -579
rect 796 -599 797 -595
rect 799 -583 800 -579
rect 799 -599 804 -583
rect 822 -595 827 -579
rect 826 -599 827 -595
rect 829 -583 830 -579
rect 829 -599 834 -583
rect 842 -595 847 -563
rect 846 -599 847 -595
rect 849 -563 851 -559
rect 855 -563 857 -559
rect 849 -599 857 -563
rect 859 -563 860 -559
rect 859 -599 864 -563
rect 868 -595 873 -559
rect 872 -599 873 -595
rect 875 -595 883 -559
rect 875 -599 877 -595
rect 881 -599 883 -595
rect 885 -563 886 -559
rect 885 -599 890 -563
rect 447 -629 452 -613
rect 451 -633 452 -629
rect 454 -617 456 -613
rect 460 -617 462 -613
rect 454 -633 462 -617
rect 464 -629 469 -613
rect 464 -633 465 -629
rect 473 -629 478 -613
rect 477 -633 478 -629
rect 480 -617 481 -613
rect 702 -606 718 -602
rect 702 -607 722 -606
rect 702 -610 722 -609
rect 480 -633 485 -617
rect 518 -618 519 -614
rect 514 -634 519 -618
rect 521 -630 526 -614
rect 632 -617 633 -613
rect 521 -634 522 -630
rect 575 -630 576 -626
rect 266 -640 286 -639
rect 270 -644 286 -640
rect 321 -640 341 -639
rect 325 -644 341 -640
rect 571 -646 576 -630
rect 578 -642 583 -626
rect 578 -646 579 -642
rect 628 -653 633 -617
rect 635 -649 643 -613
rect 635 -653 637 -649
rect 641 -653 643 -649
rect 645 -649 650 -613
rect 645 -653 646 -649
rect 658 -617 659 -613
rect 654 -653 659 -617
rect 661 -617 663 -613
rect 667 -617 669 -613
rect 661 -653 669 -617
rect 671 -617 672 -613
rect 706 -614 722 -610
rect 671 -649 676 -617
rect 671 -653 672 -649
rect 688 -637 689 -633
rect 684 -653 689 -637
rect 691 -649 696 -633
rect 691 -653 692 -649
rect 718 -637 719 -633
rect 714 -653 719 -637
rect 721 -649 726 -633
rect 721 -653 722 -649
rect 762 -637 763 -633
rect 758 -653 763 -637
rect 765 -649 770 -633
rect 765 -653 766 -649
rect 408 -663 409 -659
rect 404 -699 409 -663
rect 411 -699 419 -659
rect 421 -695 426 -659
rect 467 -663 468 -659
rect 463 -679 468 -663
rect 470 -675 478 -659
rect 470 -679 472 -675
rect 476 -679 478 -675
rect 480 -663 481 -659
rect 480 -679 485 -663
rect 508 -663 509 -659
rect 421 -699 422 -695
rect 436 -683 437 -679
rect 432 -699 437 -683
rect 439 -695 444 -679
rect 439 -699 440 -695
rect 504 -699 509 -663
rect 511 -699 519 -659
rect 521 -695 526 -659
rect 521 -699 522 -695
rect 536 -683 537 -679
rect 532 -699 537 -683
rect 539 -695 544 -679
rect 539 -699 540 -695
rect 575 -685 576 -681
rect 187 -729 188 -725
rect 183 -745 188 -729
rect 190 -741 195 -725
rect 190 -745 191 -741
rect 231 -729 232 -725
rect 227 -745 232 -729
rect 234 -741 239 -725
rect 234 -745 235 -741
rect 261 -729 262 -725
rect 257 -745 262 -729
rect 264 -741 269 -725
rect 264 -745 265 -741
rect 281 -729 282 -725
rect 277 -761 282 -729
rect 231 -768 247 -764
rect 281 -765 282 -761
rect 284 -761 292 -725
rect 284 -765 286 -761
rect 290 -765 292 -761
rect 294 -761 299 -725
rect 294 -765 295 -761
rect 307 -729 308 -725
rect 303 -765 308 -729
rect 310 -729 312 -725
rect 316 -729 318 -725
rect 310 -765 318 -729
rect 320 -761 325 -725
rect 571 -701 576 -685
rect 578 -697 583 -681
rect 578 -701 579 -697
rect 590 -697 595 -681
rect 594 -701 595 -697
rect 597 -697 602 -681
rect 597 -701 598 -697
rect 343 -755 379 -751
rect 343 -756 383 -755
rect 463 -755 479 -751
rect 463 -756 483 -755
rect 320 -765 321 -761
rect 343 -766 383 -758
rect 463 -760 483 -758
rect 467 -764 483 -760
rect 463 -766 483 -764
rect 231 -769 251 -768
rect 343 -769 383 -768
rect 231 -772 251 -771
rect 235 -776 251 -772
rect 343 -773 379 -769
rect 463 -769 483 -768
rect 463 -773 479 -769
rect 300 -789 316 -785
rect 300 -790 320 -789
rect 300 -793 320 -792
rect 304 -797 320 -793
rect 360 -832 376 -828
rect 498 -832 514 -828
rect 356 -833 376 -832
rect 356 -836 376 -835
rect 356 -840 372 -836
rect 395 -848 400 -832
rect 399 -852 400 -848
rect 402 -836 403 -832
rect 402 -852 407 -836
rect 471 -836 472 -832
rect 467 -852 472 -836
rect 474 -848 479 -832
rect 498 -833 518 -832
rect 498 -836 518 -835
rect 502 -840 518 -836
rect 474 -852 475 -848
rect 360 -862 376 -858
rect 356 -863 376 -862
rect 498 -862 514 -858
rect 498 -863 518 -862
rect 356 -866 376 -865
rect 356 -870 372 -866
rect 498 -866 518 -865
rect 502 -870 518 -866
rect 360 -882 392 -878
rect 356 -883 396 -882
rect 356 -887 396 -885
rect 356 -891 392 -887
rect 482 -882 514 -878
rect 478 -883 518 -882
rect 478 -887 518 -885
rect 356 -893 396 -891
rect 356 -896 396 -895
rect 356 -900 392 -896
rect 482 -891 518 -887
rect 478 -893 518 -891
rect 478 -896 518 -895
rect 482 -900 518 -896
rect 360 -908 396 -904
rect 356 -909 396 -908
rect 356 -913 396 -911
rect 360 -917 396 -913
rect 356 -919 396 -917
rect 416 -917 421 -901
rect 420 -921 421 -917
rect 423 -905 424 -901
rect 423 -921 428 -905
rect 450 -905 451 -901
rect 446 -921 451 -905
rect 453 -917 458 -901
rect 478 -908 514 -904
rect 478 -909 518 -908
rect 453 -921 454 -917
rect 478 -913 518 -911
rect 478 -917 514 -913
rect 478 -919 518 -917
rect 356 -922 396 -921
rect 356 -926 392 -922
rect 478 -922 518 -921
rect 482 -926 518 -922
<< ndcontact >>
rect 293 -92 297 -88
rect 514 -92 518 -88
rect 299 -101 303 -97
rect 508 -101 512 -97
rect 293 -118 297 -114
rect 299 -127 303 -123
rect 514 -118 518 -114
rect 384 -135 388 -131
rect 392 -129 396 -125
rect 415 -129 419 -125
rect 508 -127 512 -123
rect 423 -135 427 -131
rect 292 -148 296 -144
rect 515 -148 519 -144
rect 292 -157 296 -153
rect 515 -157 519 -153
rect 308 -166 312 -162
rect 292 -178 296 -174
rect 292 -187 296 -183
rect 499 -166 503 -162
rect 515 -178 519 -174
rect 308 -196 312 -192
rect 515 -187 519 -183
rect 363 -204 367 -200
rect 371 -198 375 -194
rect 436 -198 440 -194
rect 499 -196 503 -192
rect 444 -204 448 -200
rect 248 -221 252 -217
rect 242 -229 246 -225
rect 575 -237 579 -233
rect 179 -242 183 -238
rect 584 -243 588 -239
rect 173 -250 177 -246
rect 399 -251 403 -247
rect 414 -251 418 -247
rect 420 -260 424 -256
rect 601 -237 605 -233
rect 610 -243 614 -239
rect 631 -236 635 -232
rect 640 -236 644 -232
rect 649 -252 653 -248
rect 661 -236 665 -232
rect 670 -236 674 -232
rect 679 -252 683 -248
rect 705 -246 709 -242
rect 713 -252 717 -248
rect 383 -269 387 -265
rect 414 -269 418 -265
rect 147 -305 151 -301
rect 69 -312 73 -308
rect 155 -311 159 -307
rect 181 -305 185 -301
rect 75 -320 79 -316
rect 190 -321 194 -317
rect 199 -321 203 -317
rect 211 -305 215 -301
rect 220 -321 224 -317
rect 229 -321 233 -317
rect 138 -333 142 -329
rect 144 -341 148 -337
rect 250 -314 254 -310
rect 259 -320 263 -316
rect 276 -314 280 -310
rect 285 -320 289 -316
rect 786 -265 790 -261
rect 792 -273 796 -269
rect 855 -286 859 -282
rect 687 -307 691 -303
rect 681 -315 685 -311
rect 618 -328 622 -324
rect 337 -336 341 -332
rect 355 -352 359 -348
rect 378 -347 382 -343
rect 386 -353 390 -349
rect 396 -360 400 -356
rect 405 -354 409 -350
rect 612 -336 616 -332
rect 861 -294 865 -290
rect 414 -360 418 -356
rect 662 -358 666 -354
rect 289 -371 293 -367
rect 471 -370 475 -366
rect 289 -379 293 -375
rect 749 -364 753 -360
rect 758 -358 762 -354
rect 479 -376 483 -372
rect 678 -376 682 -372
rect -107 -410 -103 -406
rect -98 -416 -94 -412
rect -81 -410 -77 -406
rect -72 -416 -68 -412
rect -51 -409 -47 -405
rect -42 -409 -38 -405
rect -33 -425 -29 -421
rect -21 -409 -17 -405
rect -12 -409 -8 -405
rect 32 -411 36 -407
rect 41 -405 45 -401
rect -3 -425 1 -421
rect 58 -411 62 -407
rect 67 -405 71 -401
rect 235 -390 239 -386
rect 289 -390 293 -386
rect 540 -380 544 -376
rect 775 -364 779 -360
rect 784 -358 788 -354
rect 805 -365 809 -361
rect 814 -365 818 -361
rect 823 -349 827 -345
rect 835 -365 839 -361
rect 844 -365 848 -361
rect 853 -349 857 -345
rect 879 -355 883 -351
rect 887 -349 891 -345
rect 534 -388 538 -384
rect 88 -412 92 -408
rect 97 -412 101 -408
rect 106 -396 110 -392
rect 118 -412 122 -408
rect 127 -412 131 -408
rect 136 -396 140 -392
rect 241 -398 245 -394
rect 295 -398 299 -394
rect 527 -398 531 -394
rect 533 -407 537 -403
rect 687 -402 691 -398
rect 527 -416 531 -412
rect 681 -411 685 -407
rect 687 -420 691 -416
rect 289 -436 293 -432
rect 5 -480 9 -476
rect 289 -444 293 -440
rect 452 -424 456 -420
rect 460 -424 464 -420
rect 471 -424 475 -420
rect 782 -425 786 -421
rect 791 -409 795 -405
rect 800 -409 804 -405
rect 812 -425 816 -421
rect 821 -409 825 -405
rect 830 -409 834 -405
rect 479 -430 483 -426
rect 235 -455 239 -451
rect 289 -455 293 -451
rect 560 -443 564 -439
rect 662 -443 666 -439
rect 851 -416 855 -412
rect 860 -410 864 -406
rect 877 -416 881 -412
rect 886 -410 890 -406
rect 554 -451 558 -447
rect 344 -458 348 -454
rect 241 -463 245 -459
rect 295 -463 299 -459
rect 552 -459 556 -455
rect 352 -464 356 -460
rect 678 -461 682 -457
rect -1 -488 3 -484
rect -64 -501 -60 -497
rect 536 -477 540 -473
rect 774 -480 778 -476
rect -70 -509 -66 -505
rect 48 -509 52 -505
rect 57 -503 61 -499
rect 93 -504 97 -500
rect 252 -504 256 -500
rect 66 -509 70 -505
rect 99 -513 103 -509
rect 674 -484 678 -480
rect 714 -484 718 -480
rect 486 -495 490 -491
rect 680 -492 684 -488
rect 246 -513 250 -509
rect 325 -512 329 -508
rect 48 -524 52 -520
rect -70 -531 -66 -527
rect -64 -539 -60 -535
rect 93 -522 97 -518
rect 333 -512 337 -508
rect 344 -512 348 -508
rect 528 -502 532 -498
rect 687 -502 691 -498
rect 780 -488 784 -484
rect 732 -500 736 -496
rect 843 -501 847 -497
rect 502 -513 506 -509
rect 534 -511 538 -507
rect 681 -511 685 -507
rect 849 -509 853 -505
rect 352 -518 356 -514
rect 252 -522 256 -518
rect 404 -523 408 -519
rect 412 -517 416 -513
rect 714 -515 718 -511
rect 528 -520 532 -516
rect 687 -520 691 -516
rect 723 -521 727 -517
rect 732 -515 736 -511
rect 100 -532 104 -528
rect 66 -540 70 -536
rect 106 -540 110 -536
rect -1 -552 3 -548
rect 5 -560 9 -556
rect 244 -547 248 -543
rect 495 -547 499 -543
rect 503 -547 507 -543
rect 514 -547 518 -543
rect 522 -541 526 -537
rect 849 -531 853 -527
rect 843 -539 847 -535
rect 102 -563 106 -559
rect 228 -565 232 -561
rect 404 -569 408 -565
rect 226 -573 230 -569
rect 413 -575 417 -571
rect 422 -569 426 -565
rect 118 -581 122 -577
rect 220 -581 224 -577
rect 447 -577 451 -573
rect 465 -593 469 -589
rect 780 -552 784 -548
rect 774 -560 778 -556
rect 665 -585 669 -581
rect -107 -630 -103 -626
rect -98 -624 -94 -620
rect -81 -630 -77 -626
rect -72 -624 -68 -620
rect 93 -604 97 -600
rect -51 -631 -47 -627
rect -42 -631 -38 -627
rect -33 -615 -29 -611
rect -21 -631 -17 -627
rect -12 -631 -8 -627
rect -3 -615 1 -611
rect 99 -613 103 -609
rect 189 -612 193 -608
rect 243 -612 247 -608
rect 93 -622 97 -618
rect 195 -620 199 -616
rect 249 -620 253 -616
rect 353 -617 357 -613
rect 353 -625 357 -621
rect 100 -632 104 -628
rect 195 -631 199 -627
rect 106 -640 110 -636
rect 195 -639 199 -635
rect 299 -636 303 -632
rect 353 -636 357 -632
rect 473 -595 477 -591
rect 481 -601 485 -597
rect 514 -601 518 -597
rect 522 -595 526 -591
rect 671 -593 675 -589
rect 734 -606 738 -602
rect 305 -644 309 -640
rect 359 -644 363 -640
rect 740 -614 744 -610
rect 782 -615 786 -611
rect 791 -631 795 -627
rect 800 -631 804 -627
rect 812 -615 816 -611
rect 821 -631 825 -627
rect 830 -631 834 -627
rect 851 -624 855 -620
rect 860 -630 864 -626
rect 877 -624 881 -620
rect 886 -630 890 -626
rect 183 -713 187 -709
rect 191 -707 195 -703
rect 217 -713 221 -709
rect 226 -697 230 -693
rect 235 -697 239 -693
rect 247 -713 251 -709
rect 256 -697 260 -693
rect 265 -697 269 -693
rect 286 -704 290 -700
rect 295 -698 299 -694
rect 312 -704 316 -700
rect 321 -698 325 -694
rect 571 -669 575 -665
rect 579 -663 583 -659
rect 209 -768 213 -764
rect 404 -728 408 -724
rect 413 -722 417 -718
rect 432 -721 436 -717
rect 440 -715 444 -711
rect 463 -719 467 -715
rect 481 -703 485 -699
rect 628 -684 632 -680
rect 637 -678 641 -674
rect 422 -728 426 -724
rect 504 -728 508 -724
rect 513 -722 517 -718
rect 532 -721 536 -717
rect 540 -715 544 -711
rect 654 -684 658 -680
rect 663 -678 667 -674
rect 684 -685 688 -681
rect 693 -685 697 -681
rect 702 -669 706 -665
rect 714 -685 718 -681
rect 723 -685 727 -681
rect 732 -669 736 -665
rect 758 -675 762 -671
rect 766 -669 770 -665
rect 522 -728 526 -724
rect 571 -723 575 -719
rect 579 -717 583 -713
rect 590 -717 594 -713
rect 598 -717 602 -713
rect 408 -755 412 -751
rect 439 -755 443 -751
rect 402 -764 406 -760
rect 215 -776 219 -772
rect 408 -773 412 -769
rect 423 -773 427 -769
rect 278 -789 282 -785
rect 284 -797 288 -793
rect 395 -814 399 -810
rect 340 -822 344 -818
rect 403 -820 407 -816
rect 467 -820 471 -816
rect 475 -814 479 -810
rect 324 -831 328 -827
rect 530 -822 534 -818
rect 324 -840 328 -836
rect 340 -852 344 -848
rect 546 -831 550 -827
rect 546 -840 550 -836
rect 530 -852 534 -848
rect 324 -861 328 -857
rect 546 -861 550 -857
rect 324 -870 328 -866
rect 546 -870 550 -866
rect 416 -883 420 -879
rect 331 -891 335 -887
rect 424 -889 428 -885
rect 446 -889 450 -885
rect 454 -883 458 -879
rect 325 -900 329 -896
rect 539 -891 543 -887
rect 545 -900 549 -896
rect 331 -917 335 -913
rect 539 -917 543 -913
rect 325 -926 329 -922
rect 545 -926 549 -922
<< pdcontact >>
rect 360 -92 364 -88
rect 447 -92 451 -88
rect 324 -101 328 -97
rect 384 -97 388 -93
rect 324 -110 328 -106
rect 392 -113 396 -109
rect 415 -113 419 -109
rect 423 -97 427 -93
rect 483 -101 487 -97
rect 483 -110 487 -106
rect 360 -118 364 -114
rect 360 -127 364 -123
rect 447 -118 451 -114
rect 324 -136 328 -132
rect 360 -136 364 -132
rect 447 -127 451 -123
rect 447 -136 451 -132
rect 483 -136 487 -132
rect 340 -148 344 -144
rect 467 -148 471 -144
rect 324 -156 328 -152
rect 483 -156 487 -152
rect 363 -166 367 -162
rect 340 -178 344 -174
rect 371 -182 375 -178
rect 436 -182 440 -178
rect 444 -166 448 -162
rect 467 -178 471 -174
rect 324 -186 328 -182
rect 483 -186 487 -182
rect 264 -221 268 -217
rect 280 -229 284 -225
rect 195 -242 199 -238
rect 211 -250 215 -246
rect 241 -253 245 -249
rect 147 -289 151 -285
rect 155 -273 159 -269
rect 191 -289 195 -285
rect 199 -273 203 -269
rect 221 -289 225 -285
rect 229 -273 233 -269
rect 241 -289 245 -285
rect 250 -253 254 -249
rect 259 -253 263 -249
rect 267 -289 271 -285
rect 276 -289 280 -285
rect 285 -253 289 -249
rect 343 -251 347 -247
rect 479 -251 483 -247
rect 359 -260 363 -256
rect 343 -269 347 -265
rect 443 -269 447 -265
rect 53 -312 57 -308
rect 37 -320 41 -316
rect 122 -333 126 -329
rect 32 -344 36 -340
rect 41 -380 45 -376
rect 50 -380 54 -376
rect 58 -344 62 -340
rect 67 -344 71 -340
rect 76 -344 80 -340
rect 106 -341 110 -337
rect 337 -296 341 -292
rect 346 -312 350 -308
rect 355 -296 359 -292
rect 378 -331 382 -327
rect 386 -315 390 -311
rect 396 -331 400 -327
rect 414 -295 418 -291
rect 575 -304 579 -300
rect 584 -268 588 -264
rect 593 -268 597 -264
rect 601 -304 605 -300
rect 610 -304 614 -300
rect 619 -268 623 -264
rect 631 -284 635 -280
rect 639 -268 643 -264
rect 661 -284 665 -280
rect 669 -268 673 -264
rect 705 -284 709 -280
rect 713 -268 717 -264
rect 770 -265 774 -261
rect 754 -273 758 -269
rect 839 -286 843 -282
rect 619 -304 623 -300
rect 749 -297 753 -293
rect 649 -307 653 -303
rect 665 -315 669 -311
rect 580 -328 584 -324
rect 471 -353 475 -349
rect 479 -337 483 -333
rect 596 -336 600 -332
rect 758 -333 762 -329
rect 767 -333 771 -329
rect 775 -297 779 -293
rect 784 -297 788 -293
rect 793 -297 797 -293
rect 823 -294 827 -290
rect 793 -333 797 -329
rect 805 -317 809 -313
rect 813 -333 817 -329
rect 835 -317 839 -313
rect 843 -333 847 -329
rect 879 -317 883 -313
rect 887 -333 891 -329
rect 76 -380 80 -376
rect 88 -364 92 -360
rect 96 -380 100 -376
rect 118 -364 122 -360
rect 622 -358 626 -354
rect 273 -371 277 -367
rect 126 -380 130 -376
rect 273 -379 277 -375
rect 638 -367 642 -363
rect 622 -376 626 -372
rect 218 -390 222 -386
rect 273 -390 277 -386
rect 556 -380 560 -376
rect 572 -388 576 -384
rect 202 -398 206 -394
rect 257 -398 261 -394
rect 452 -408 456 -404
rect 460 -408 464 -404
rect 471 -408 475 -404
rect 479 -392 483 -388
rect 556 -398 560 -394
rect 658 -402 662 -398
rect 592 -416 596 -412
rect 622 -420 626 -416
rect 273 -436 277 -432
rect -107 -477 -103 -473
rect -98 -441 -94 -437
rect -89 -441 -85 -437
rect -81 -477 -77 -473
rect -72 -477 -68 -473
rect -63 -441 -59 -437
rect -51 -457 -47 -453
rect -43 -441 -39 -437
rect -21 -457 -17 -453
rect -13 -441 -9 -437
rect -63 -477 -59 -473
rect -33 -480 -29 -476
rect 48 -480 52 -476
rect 273 -444 277 -440
rect 344 -441 348 -437
rect 352 -425 356 -421
rect 218 -455 222 -451
rect 273 -455 277 -451
rect 576 -443 580 -439
rect 622 -443 626 -439
rect 714 -444 718 -440
rect 592 -451 596 -447
rect 638 -452 642 -448
rect 202 -463 206 -459
rect 257 -463 261 -459
rect 592 -459 596 -455
rect 622 -461 626 -457
rect 723 -460 727 -456
rect 732 -444 736 -440
rect 792 -441 796 -437
rect 800 -457 804 -453
rect 822 -441 826 -437
rect 830 -457 834 -453
rect 842 -441 846 -437
rect 576 -468 580 -464
rect 66 -480 70 -476
rect -17 -488 -13 -484
rect -102 -501 -98 -497
rect 325 -496 329 -492
rect 333 -496 337 -492
rect 344 -496 348 -492
rect 352 -480 356 -476
rect 592 -477 596 -473
rect 404 -485 408 -481
rect -86 -509 -82 -505
rect 158 -504 162 -500
rect 187 -504 191 -500
rect 658 -484 662 -480
rect 446 -495 450 -491
rect 642 -492 646 -488
rect 412 -501 416 -497
rect -86 -531 -82 -527
rect -102 -539 -98 -535
rect 122 -522 126 -518
rect 223 -522 227 -518
rect 462 -504 466 -500
rect 557 -502 561 -498
rect 658 -502 662 -498
rect 812 -480 816 -476
rect 842 -477 846 -473
rect 851 -477 855 -473
rect 860 -477 864 -473
rect 868 -441 872 -437
rect 877 -441 881 -437
rect 886 -477 890 -473
rect 796 -488 800 -484
rect 881 -501 885 -497
rect 446 -513 450 -509
rect 865 -509 869 -505
rect 571 -520 575 -516
rect 593 -520 597 -516
rect 622 -520 626 -516
rect 138 -532 142 -528
rect 122 -540 126 -536
rect -17 -552 -13 -548
rect -107 -563 -103 -559
rect -98 -599 -94 -595
rect -89 -599 -85 -595
rect -81 -563 -77 -559
rect -72 -563 -68 -559
rect -63 -563 -59 -559
rect -33 -560 -29 -556
rect 188 -547 192 -543
rect 865 -531 869 -527
rect 881 -539 885 -535
rect 714 -544 718 -540
rect 204 -556 208 -552
rect -63 -599 -59 -595
rect -51 -583 -47 -579
rect -43 -599 -39 -595
rect -21 -583 -17 -579
rect 48 -580 52 -576
rect 57 -564 61 -560
rect 158 -563 162 -559
rect 188 -565 192 -561
rect 495 -563 499 -559
rect 142 -572 146 -568
rect 188 -573 192 -569
rect 66 -580 70 -576
rect 158 -581 162 -577
rect 204 -581 208 -577
rect 503 -563 507 -559
rect 514 -563 518 -559
rect 522 -579 526 -575
rect 732 -544 736 -540
rect 796 -552 800 -548
rect 812 -560 816 -556
rect 842 -563 846 -559
rect 649 -585 653 -581
rect -13 -599 -9 -595
rect 158 -604 162 -600
rect 227 -612 231 -608
rect 282 -612 286 -608
rect 122 -622 126 -618
rect 211 -620 215 -616
rect 266 -620 270 -616
rect 337 -617 341 -613
rect 337 -625 341 -621
rect 138 -632 142 -628
rect 211 -631 215 -627
rect 122 -640 126 -636
rect 211 -639 215 -635
rect 282 -636 286 -632
rect 337 -636 341 -632
rect 404 -634 408 -630
rect 422 -598 426 -594
rect 633 -593 637 -589
rect 792 -599 796 -595
rect 800 -583 804 -579
rect 822 -599 826 -595
rect 830 -583 834 -579
rect 842 -599 846 -595
rect 851 -563 855 -559
rect 860 -563 864 -559
rect 868 -599 872 -595
rect 877 -599 881 -595
rect 886 -563 890 -559
rect 447 -633 451 -629
rect 456 -617 460 -613
rect 465 -633 469 -629
rect 473 -633 477 -629
rect 481 -617 485 -613
rect 718 -606 722 -602
rect 514 -618 518 -614
rect 628 -617 632 -613
rect 522 -634 526 -630
rect 571 -630 575 -626
rect 266 -644 270 -640
rect 321 -644 325 -640
rect 579 -646 583 -642
rect 637 -653 641 -649
rect 646 -653 650 -649
rect 654 -617 658 -613
rect 663 -617 667 -613
rect 672 -617 676 -613
rect 702 -614 706 -610
rect 672 -653 676 -649
rect 684 -637 688 -633
rect 692 -653 696 -649
rect 714 -637 718 -633
rect 722 -653 726 -649
rect 758 -637 762 -633
rect 766 -653 770 -649
rect 404 -663 408 -659
rect 463 -663 467 -659
rect 472 -679 476 -675
rect 481 -663 485 -659
rect 504 -663 508 -659
rect 422 -699 426 -695
rect 432 -683 436 -679
rect 440 -699 444 -695
rect 522 -699 526 -695
rect 532 -683 536 -679
rect 540 -699 544 -695
rect 571 -685 575 -681
rect 183 -729 187 -725
rect 191 -745 195 -741
rect 227 -729 231 -725
rect 235 -745 239 -741
rect 257 -729 261 -725
rect 265 -745 269 -741
rect 277 -729 281 -725
rect 247 -768 251 -764
rect 277 -765 281 -761
rect 286 -765 290 -761
rect 295 -765 299 -761
rect 303 -729 307 -725
rect 312 -729 316 -725
rect 579 -701 583 -697
rect 590 -701 594 -697
rect 598 -701 602 -697
rect 379 -755 383 -751
rect 479 -755 483 -751
rect 321 -765 325 -761
rect 463 -764 467 -760
rect 231 -776 235 -772
rect 379 -773 383 -769
rect 479 -773 483 -769
rect 316 -789 320 -785
rect 300 -797 304 -793
rect 356 -832 360 -828
rect 514 -832 518 -828
rect 372 -840 376 -836
rect 395 -852 399 -848
rect 403 -836 407 -832
rect 467 -836 471 -832
rect 498 -840 502 -836
rect 475 -852 479 -848
rect 356 -862 360 -858
rect 514 -862 518 -858
rect 372 -870 376 -866
rect 498 -870 502 -866
rect 356 -882 360 -878
rect 392 -882 396 -878
rect 392 -891 396 -887
rect 478 -882 482 -878
rect 514 -882 518 -878
rect 392 -900 396 -896
rect 478 -891 482 -887
rect 478 -900 482 -896
rect 356 -908 360 -904
rect 356 -917 360 -913
rect 416 -921 420 -917
rect 424 -905 428 -901
rect 446 -905 450 -901
rect 514 -908 518 -904
rect 454 -921 458 -917
rect 514 -917 518 -913
rect 392 -926 396 -922
rect 478 -926 482 -922
<< polysilicon >>
rect 389 -93 391 -89
rect 420 -93 422 -89
rect 290 -95 293 -93
rect 303 -95 324 -93
rect 364 -95 367 -93
rect 275 -105 324 -103
rect 364 -105 367 -103
rect 444 -95 447 -93
rect 487 -95 508 -93
rect 518 -95 521 -93
rect 444 -105 447 -103
rect 487 -105 536 -103
rect 290 -121 293 -119
rect 303 -121 324 -119
rect 364 -121 367 -119
rect 389 -125 391 -113
rect 420 -125 422 -113
rect 444 -121 447 -119
rect 487 -121 508 -119
rect 518 -121 521 -119
rect 275 -131 324 -129
rect 364 -131 367 -129
rect 444 -131 447 -129
rect 487 -131 536 -129
rect 389 -139 391 -135
rect 420 -139 422 -135
rect 289 -151 292 -149
rect 312 -151 324 -149
rect 344 -151 348 -149
rect 463 -151 467 -149
rect 487 -151 499 -149
rect 519 -151 522 -149
rect 275 -161 292 -159
rect 312 -161 315 -159
rect 368 -162 370 -158
rect 441 -162 443 -158
rect 496 -161 499 -159
rect 519 -161 536 -159
rect 289 -181 292 -179
rect 312 -181 324 -179
rect 344 -181 348 -179
rect 463 -181 467 -179
rect 487 -181 499 -179
rect 519 -181 522 -179
rect 275 -191 292 -189
rect 312 -191 315 -189
rect 368 -194 370 -182
rect 441 -194 443 -182
rect 496 -191 499 -189
rect 519 -191 536 -189
rect 368 -208 370 -204
rect 441 -208 443 -204
rect 238 -224 242 -222
rect 252 -224 264 -222
rect 284 -224 288 -222
rect 580 -233 582 -230
rect 169 -245 173 -243
rect 183 -245 195 -243
rect 215 -245 219 -243
rect 246 -249 248 -246
rect 256 -249 258 -246
rect 272 -249 274 -246
rect 282 -249 284 -246
rect 152 -269 154 -265
rect 196 -269 198 -265
rect 226 -269 228 -265
rect 339 -254 343 -252
rect 363 -254 383 -252
rect 403 -254 406 -252
rect 411 -254 414 -252
rect 424 -254 443 -252
rect 483 -254 486 -252
rect 339 -264 343 -262
rect 363 -264 383 -262
rect 403 -264 406 -262
rect 411 -264 414 -262
rect 424 -264 443 -262
rect 483 -264 486 -262
rect 580 -264 582 -243
rect 590 -264 592 -215
rect 606 -233 608 -230
rect 606 -264 608 -243
rect 616 -264 618 -215
rect 636 -232 638 -229
rect 646 -232 648 -215
rect 666 -232 668 -229
rect 676 -232 678 -215
rect 710 -242 712 -238
rect 636 -264 638 -252
rect 646 -255 648 -252
rect 666 -264 668 -252
rect 676 -255 678 -252
rect 710 -264 712 -252
rect 152 -301 154 -289
rect 186 -301 188 -298
rect 196 -301 198 -289
rect 216 -301 218 -298
rect 226 -301 228 -289
rect 33 -315 37 -313
rect 57 -315 69 -313
rect 79 -315 83 -313
rect 152 -315 154 -311
rect 102 -336 106 -334
rect 126 -336 138 -334
rect 148 -336 152 -334
rect 37 -340 39 -337
rect 47 -340 49 -337
rect 63 -340 65 -337
rect 73 -340 75 -337
rect 186 -338 188 -321
rect 196 -324 198 -321
rect 216 -338 218 -321
rect 226 -324 228 -321
rect 246 -338 248 -289
rect 256 -310 258 -289
rect 256 -323 258 -320
rect 272 -338 274 -289
rect 282 -310 284 -289
rect 342 -292 344 -288
rect 352 -292 354 -288
rect 401 -291 403 -288
rect 411 -291 413 -288
rect 383 -311 385 -307
rect 282 -323 284 -320
rect 342 -332 344 -312
rect 352 -332 354 -312
rect 750 -268 754 -266
rect 774 -268 786 -266
rect 796 -268 800 -266
rect 636 -288 638 -284
rect 666 -288 668 -284
rect 710 -288 712 -284
rect 819 -289 823 -287
rect 843 -289 855 -287
rect 865 -289 869 -287
rect 754 -293 756 -290
rect 764 -293 766 -290
rect 780 -293 782 -290
rect 790 -293 792 -290
rect 580 -307 582 -304
rect 590 -307 592 -304
rect 606 -307 608 -304
rect 616 -307 618 -304
rect 645 -310 649 -308
rect 669 -310 681 -308
rect 691 -310 695 -308
rect 383 -343 385 -331
rect 342 -355 344 -352
rect 352 -355 354 -352
rect 401 -350 403 -331
rect 411 -350 413 -331
rect 476 -333 478 -329
rect 576 -331 580 -329
rect 600 -331 612 -329
rect 622 -331 626 -329
rect 93 -360 95 -356
rect 123 -360 125 -356
rect 383 -357 385 -353
rect 810 -313 812 -309
rect 840 -313 842 -309
rect 884 -313 886 -309
rect 401 -363 403 -360
rect 411 -363 413 -360
rect 476 -366 478 -353
rect 754 -354 756 -333
rect 618 -361 622 -359
rect 642 -361 662 -359
rect 682 -361 685 -359
rect 245 -374 257 -372
rect 277 -374 280 -372
rect 286 -374 289 -372
rect 299 -374 305 -372
rect 754 -367 756 -364
rect 618 -371 622 -369
rect 642 -371 662 -369
rect 682 -371 685 -369
rect -102 -406 -100 -403
rect -102 -437 -100 -416
rect -92 -437 -90 -388
rect -76 -406 -74 -403
rect -76 -437 -74 -416
rect -66 -437 -64 -388
rect -46 -405 -44 -402
rect -36 -405 -34 -388
rect -16 -405 -14 -402
rect -6 -405 -4 -388
rect 37 -401 39 -380
rect 37 -414 39 -411
rect -46 -437 -44 -425
rect -36 -428 -34 -425
rect -16 -437 -14 -425
rect -6 -428 -4 -425
rect 47 -429 49 -380
rect 63 -401 65 -380
rect 63 -414 65 -411
rect 73 -429 75 -380
rect 93 -392 95 -380
rect 103 -392 105 -389
rect 123 -392 125 -380
rect 133 -392 135 -389
rect 457 -388 459 -376
rect 476 -380 478 -376
rect 530 -383 534 -381
rect 544 -383 556 -381
rect 576 -383 580 -381
rect 764 -382 766 -333
rect 780 -354 782 -333
rect 780 -367 782 -364
rect 790 -382 792 -333
rect 810 -345 812 -333
rect 820 -345 822 -342
rect 840 -345 842 -333
rect 850 -345 852 -342
rect 884 -345 886 -333
rect 884 -359 886 -355
rect 810 -368 812 -365
rect 820 -382 822 -365
rect 840 -368 842 -365
rect 850 -382 852 -365
rect 476 -388 478 -384
rect 198 -393 202 -391
rect 222 -393 235 -391
rect 245 -393 249 -391
rect 253 -393 257 -391
rect 277 -393 289 -391
rect 299 -393 302 -391
rect 524 -401 527 -399
rect 537 -401 556 -399
rect 596 -401 599 -399
rect 457 -411 459 -408
rect 93 -415 95 -412
rect 103 -429 105 -412
rect 123 -415 125 -412
rect 133 -429 135 -412
rect 349 -421 351 -417
rect 457 -420 459 -417
rect 476 -420 478 -408
rect 619 -405 622 -403
rect 662 -405 681 -403
rect 691 -405 694 -403
rect 787 -405 789 -388
rect 797 -405 799 -402
rect 817 -405 819 -388
rect 827 -405 829 -402
rect 524 -411 527 -409
rect 537 -411 556 -409
rect 596 -411 599 -409
rect 619 -415 622 -413
rect 662 -415 681 -413
rect 691 -415 694 -413
rect 53 -440 55 -437
rect 63 -440 65 -437
rect 245 -439 257 -437
rect 277 -439 280 -437
rect 286 -439 289 -437
rect 299 -439 305 -437
rect -46 -461 -44 -457
rect -16 -461 -14 -457
rect -102 -480 -100 -477
rect -92 -480 -90 -477
rect -76 -480 -74 -477
rect -66 -480 -64 -477
rect 787 -428 789 -425
rect 457 -436 459 -430
rect 476 -433 478 -430
rect 349 -454 351 -441
rect 719 -440 721 -436
rect 729 -440 731 -436
rect 797 -437 799 -425
rect 817 -428 819 -425
rect 827 -437 829 -425
rect 847 -437 849 -388
rect 857 -406 859 -403
rect 857 -437 859 -416
rect 873 -437 875 -388
rect 883 -406 885 -403
rect 883 -437 885 -416
rect 550 -446 554 -444
rect 564 -446 576 -444
rect 596 -446 600 -444
rect 618 -446 622 -444
rect 642 -446 662 -444
rect 682 -446 685 -444
rect 198 -458 202 -456
rect 222 -458 235 -456
rect 245 -458 249 -456
rect 253 -458 257 -456
rect 277 -458 289 -456
rect 299 -458 302 -456
rect 618 -456 622 -454
rect 642 -456 662 -454
rect 682 -456 685 -454
rect 533 -462 536 -460
rect 556 -462 576 -460
rect 596 -462 600 -460
rect 330 -476 332 -464
rect 349 -468 351 -464
rect 533 -472 536 -470
rect 556 -472 576 -470
rect 596 -472 600 -470
rect 349 -476 351 -472
rect -37 -483 -33 -481
rect -13 -483 -1 -481
rect 9 -483 13 -481
rect 53 -499 55 -480
rect 63 -499 65 -480
rect 409 -481 411 -477
rect 719 -480 721 -460
rect 729 -480 731 -460
rect 797 -461 799 -457
rect 827 -461 829 -457
rect 330 -499 332 -496
rect -106 -504 -102 -502
rect -82 -504 -70 -502
rect -60 -504 -56 -502
rect 90 -507 93 -505
rect 103 -507 122 -505
rect 162 -507 165 -505
rect 184 -507 187 -505
rect 227 -507 246 -505
rect 256 -507 259 -505
rect 53 -512 55 -509
rect 63 -512 65 -509
rect 330 -508 332 -505
rect 349 -508 351 -496
rect 638 -487 642 -485
rect 662 -487 674 -485
rect 684 -487 688 -485
rect 442 -498 446 -496
rect 466 -498 486 -496
rect 506 -498 509 -496
rect 90 -517 93 -515
rect 103 -517 122 -515
rect 162 -517 165 -515
rect 184 -517 187 -515
rect 227 -517 246 -515
rect 256 -517 259 -515
rect 53 -520 55 -517
rect 63 -520 65 -517
rect -106 -534 -102 -532
rect -82 -534 -70 -532
rect -60 -534 -56 -532
rect 409 -513 411 -501
rect 847 -480 849 -477
rect 857 -480 859 -477
rect 873 -480 875 -477
rect 883 -480 885 -477
rect 770 -483 774 -481
rect 784 -483 796 -481
rect 816 -483 820 -481
rect 719 -503 721 -500
rect 729 -503 731 -500
rect 525 -505 528 -503
rect 538 -505 557 -503
rect 597 -505 600 -503
rect 619 -505 622 -503
rect 662 -505 681 -503
rect 691 -505 694 -503
rect 839 -504 843 -502
rect 853 -504 865 -502
rect 885 -504 889 -502
rect 442 -508 446 -506
rect 466 -508 486 -506
rect 506 -508 509 -506
rect 719 -511 721 -508
rect 729 -511 731 -508
rect 330 -524 332 -518
rect 349 -521 351 -518
rect 525 -515 528 -513
rect 538 -515 557 -513
rect 597 -515 600 -513
rect 619 -515 622 -513
rect 662 -515 681 -513
rect 691 -515 694 -513
rect 409 -527 411 -523
rect 96 -535 100 -533
rect 110 -535 122 -533
rect 142 -535 146 -533
rect 500 -537 502 -531
rect 519 -537 521 -534
rect -37 -555 -33 -553
rect -13 -555 -1 -553
rect 9 -555 13 -553
rect -102 -559 -100 -556
rect -92 -559 -90 -556
rect -76 -559 -74 -556
rect -66 -559 -64 -556
rect 53 -560 55 -540
rect 63 -560 65 -540
rect 719 -540 721 -521
rect 729 -540 731 -521
rect 839 -534 843 -532
rect 853 -534 865 -532
rect 885 -534 889 -532
rect 184 -550 188 -548
rect 208 -550 228 -548
rect 248 -550 251 -548
rect 500 -550 502 -547
rect -46 -579 -44 -575
rect -16 -579 -14 -575
rect 184 -560 188 -558
rect 208 -560 228 -558
rect 248 -560 251 -558
rect 500 -559 502 -556
rect 519 -559 521 -547
rect 99 -566 102 -564
rect 122 -566 142 -564
rect 162 -566 166 -564
rect 409 -565 411 -562
rect 419 -565 421 -562
rect 99 -576 102 -574
rect 122 -576 142 -574
rect 162 -576 166 -574
rect 184 -576 188 -574
rect 208 -576 220 -574
rect 230 -576 234 -574
rect 452 -573 454 -570
rect 462 -573 464 -570
rect 53 -584 55 -580
rect 63 -584 65 -580
rect 409 -594 411 -575
rect 419 -594 421 -575
rect 478 -591 480 -587
rect 500 -591 502 -579
rect 519 -583 521 -579
rect 770 -555 774 -553
rect 784 -555 796 -553
rect 816 -555 820 -553
rect 847 -559 849 -556
rect 857 -559 859 -556
rect 873 -559 875 -556
rect 883 -559 885 -556
rect 797 -579 799 -575
rect 827 -579 829 -575
rect 719 -583 721 -580
rect 729 -583 731 -580
rect 519 -591 521 -587
rect 629 -588 633 -586
rect 653 -588 665 -586
rect 675 -588 679 -586
rect -102 -620 -100 -599
rect -102 -633 -100 -630
rect -92 -648 -90 -599
rect -76 -620 -74 -599
rect -76 -633 -74 -630
rect -66 -648 -64 -599
rect -46 -611 -44 -599
rect -36 -611 -34 -608
rect -16 -611 -14 -599
rect 90 -607 93 -605
rect 103 -607 122 -605
rect 162 -607 165 -605
rect -6 -611 -4 -608
rect 186 -615 189 -613
rect 199 -615 211 -613
rect 231 -615 235 -613
rect 239 -615 243 -613
rect 253 -615 266 -613
rect 286 -615 290 -613
rect 90 -617 93 -615
rect 103 -617 122 -615
rect 162 -617 165 -615
rect 309 -620 321 -618
rect 341 -620 344 -618
rect 350 -620 353 -618
rect 363 -620 369 -618
rect -46 -634 -44 -631
rect -36 -648 -34 -631
rect -16 -634 -14 -631
rect -6 -648 -4 -631
rect 96 -635 100 -633
rect 110 -635 122 -633
rect 142 -635 146 -633
rect 183 -634 189 -632
rect 199 -634 202 -632
rect 208 -634 211 -632
rect 231 -634 243 -632
rect 452 -613 454 -593
rect 462 -613 464 -593
rect 478 -613 480 -601
rect 519 -614 521 -601
rect 698 -609 702 -607
rect 722 -609 734 -607
rect 744 -609 748 -607
rect 633 -613 635 -610
rect 643 -613 645 -610
rect 659 -613 661 -610
rect 669 -613 671 -610
rect 409 -637 411 -634
rect 419 -637 421 -634
rect 452 -637 454 -633
rect 462 -637 464 -633
rect 478 -637 480 -633
rect 576 -626 578 -622
rect 262 -639 266 -637
rect 286 -639 299 -637
rect 309 -639 313 -637
rect 317 -639 321 -637
rect 341 -639 353 -637
rect 363 -639 366 -637
rect 519 -638 521 -634
rect 409 -659 411 -656
rect 419 -659 421 -656
rect 468 -659 470 -655
rect 478 -659 480 -655
rect 509 -659 511 -656
rect 519 -659 521 -656
rect 576 -659 578 -646
rect 787 -611 789 -608
rect 797 -611 799 -599
rect 817 -611 819 -608
rect 827 -611 829 -599
rect 689 -633 691 -629
rect 719 -633 721 -629
rect 763 -633 765 -629
rect 787 -648 789 -631
rect 797 -634 799 -631
rect 817 -648 819 -631
rect 827 -634 829 -631
rect 847 -648 849 -599
rect 857 -620 859 -599
rect 857 -633 859 -630
rect 873 -648 875 -599
rect 883 -620 885 -599
rect 883 -633 885 -630
rect 222 -693 224 -676
rect 232 -693 234 -690
rect 252 -693 254 -676
rect 262 -693 264 -690
rect 188 -703 190 -699
rect 188 -725 190 -713
rect 222 -716 224 -713
rect 232 -725 234 -713
rect 252 -716 254 -713
rect 262 -725 264 -713
rect 282 -725 284 -676
rect 292 -694 294 -691
rect 292 -725 294 -704
rect 308 -725 310 -676
rect 318 -694 320 -691
rect 437 -679 439 -675
rect 468 -699 470 -679
rect 478 -699 480 -679
rect 576 -673 578 -669
rect 537 -679 539 -675
rect 576 -681 578 -677
rect 595 -681 597 -669
rect 633 -674 635 -653
rect 318 -725 320 -704
rect 409 -718 411 -699
rect 419 -718 421 -699
rect 437 -711 439 -699
rect 188 -749 190 -745
rect 232 -749 234 -745
rect 262 -749 264 -745
rect 509 -718 511 -699
rect 519 -718 521 -699
rect 537 -711 539 -699
rect 633 -687 635 -684
rect 437 -725 439 -721
rect 468 -722 470 -719
rect 478 -722 480 -719
rect 576 -713 578 -701
rect 595 -704 597 -701
rect 643 -702 645 -653
rect 659 -674 661 -653
rect 659 -687 661 -684
rect 669 -702 671 -653
rect 689 -665 691 -653
rect 699 -665 701 -662
rect 719 -665 721 -653
rect 729 -665 731 -662
rect 763 -665 765 -653
rect 763 -679 765 -675
rect 689 -688 691 -685
rect 699 -702 701 -685
rect 719 -688 721 -685
rect 729 -702 731 -685
rect 595 -713 597 -710
rect 537 -725 539 -721
rect 576 -726 578 -723
rect 409 -731 411 -728
rect 419 -731 421 -728
rect 509 -731 511 -728
rect 519 -731 521 -728
rect 595 -729 597 -723
rect 340 -758 343 -756
rect 383 -758 402 -756
rect 412 -758 415 -756
rect 420 -758 423 -756
rect 443 -758 463 -756
rect 483 -758 487 -756
rect 282 -768 284 -765
rect 292 -768 294 -765
rect 308 -768 310 -765
rect 318 -768 320 -765
rect 340 -768 343 -766
rect 383 -768 402 -766
rect 412 -768 415 -766
rect 420 -768 423 -766
rect 443 -768 463 -766
rect 483 -768 487 -766
rect 205 -771 209 -769
rect 219 -771 231 -769
rect 251 -771 255 -769
rect 274 -792 278 -790
rect 288 -792 300 -790
rect 320 -792 324 -790
rect 400 -810 402 -806
rect 472 -810 474 -806
rect 307 -825 324 -823
rect 344 -825 347 -823
rect 400 -832 402 -820
rect 472 -832 474 -820
rect 527 -825 530 -823
rect 550 -825 567 -823
rect 321 -835 324 -833
rect 344 -835 356 -833
rect 376 -835 380 -833
rect 494 -835 498 -833
rect 518 -835 530 -833
rect 550 -835 553 -833
rect 307 -855 324 -853
rect 344 -855 347 -853
rect 400 -856 402 -852
rect 472 -856 474 -852
rect 527 -855 530 -853
rect 550 -855 567 -853
rect 321 -865 324 -863
rect 344 -865 356 -863
rect 376 -865 380 -863
rect 494 -865 498 -863
rect 518 -865 530 -863
rect 550 -865 553 -863
rect 421 -879 423 -875
rect 451 -879 453 -875
rect 307 -885 356 -883
rect 396 -885 399 -883
rect 475 -885 478 -883
rect 518 -885 567 -883
rect 322 -895 325 -893
rect 335 -895 356 -893
rect 396 -895 399 -893
rect 421 -901 423 -889
rect 451 -901 453 -889
rect 475 -895 478 -893
rect 518 -895 539 -893
rect 549 -895 552 -893
rect 307 -911 356 -909
rect 396 -911 399 -909
rect 322 -921 325 -919
rect 335 -921 356 -919
rect 396 -921 399 -919
rect 475 -911 478 -909
rect 518 -911 567 -909
rect 475 -921 478 -919
rect 518 -921 539 -919
rect 549 -921 552 -919
rect 421 -925 423 -921
rect 451 -925 453 -921
<< polycontact >>
rect 307 -93 311 -89
rect 500 -93 504 -89
rect 278 -103 282 -99
rect 529 -103 533 -99
rect 308 -119 312 -115
rect 278 -129 282 -125
rect 385 -124 389 -120
rect 499 -119 503 -115
rect 422 -124 426 -120
rect 529 -129 533 -125
rect 313 -149 317 -145
rect 494 -149 498 -145
rect 278 -159 282 -155
rect 529 -159 533 -155
rect 313 -179 317 -175
rect 278 -189 282 -185
rect 494 -179 498 -175
rect 364 -193 368 -189
rect 529 -189 533 -185
rect 443 -193 447 -189
rect 586 -222 590 -218
rect 253 -228 257 -224
rect 184 -249 188 -245
rect 370 -252 374 -248
rect 425 -252 429 -248
rect 576 -251 580 -247
rect 378 -262 382 -258
rect 432 -262 436 -258
rect 612 -222 616 -218
rect 602 -252 606 -248
rect 642 -222 646 -218
rect 672 -222 676 -218
rect 632 -257 636 -253
rect 662 -257 666 -253
rect 706 -257 710 -253
rect 154 -300 158 -296
rect 198 -300 202 -296
rect 228 -300 232 -296
rect 64 -319 68 -315
rect 133 -340 137 -336
rect 188 -335 192 -331
rect 218 -335 222 -331
rect 258 -305 262 -301
rect 248 -335 252 -331
rect 284 -306 288 -302
rect 274 -335 278 -331
rect 344 -331 348 -327
rect 354 -323 358 -319
rect 781 -272 785 -268
rect 676 -308 680 -304
rect 607 -329 611 -325
rect 385 -342 389 -338
rect 403 -342 407 -338
rect 413 -349 417 -345
rect 850 -293 854 -289
rect 750 -350 754 -346
rect 478 -365 482 -361
rect 300 -372 304 -368
rect 246 -378 250 -374
rect 657 -365 661 -361
rect 649 -375 653 -371
rect -96 -395 -92 -391
rect -106 -424 -102 -420
rect -70 -395 -66 -391
rect -80 -425 -76 -421
rect -40 -395 -36 -391
rect -10 -395 -6 -391
rect 33 -397 37 -393
rect -50 -430 -46 -426
rect -20 -430 -16 -426
rect 43 -426 47 -422
rect 59 -396 63 -392
rect 69 -426 73 -422
rect 89 -391 93 -387
rect 119 -391 123 -387
rect 459 -381 463 -377
rect 760 -379 764 -375
rect 776 -349 780 -345
rect 786 -379 790 -375
rect 806 -344 810 -340
rect 836 -344 840 -340
rect 880 -344 884 -340
rect 816 -379 820 -375
rect 846 -379 850 -375
rect 545 -387 549 -383
rect 230 -397 234 -393
rect 284 -397 288 -393
rect 545 -405 549 -401
rect 99 -426 103 -422
rect 129 -426 133 -422
rect 789 -395 793 -391
rect 819 -395 823 -391
rect 478 -419 482 -415
rect 538 -415 542 -411
rect 669 -409 673 -405
rect 676 -419 680 -415
rect 300 -437 304 -433
rect -6 -481 -2 -477
rect 246 -443 250 -439
rect 453 -435 457 -431
rect 799 -430 803 -426
rect 829 -430 833 -426
rect 849 -395 853 -391
rect 859 -425 863 -421
rect 875 -395 879 -391
rect 885 -424 889 -420
rect 351 -453 355 -449
rect 565 -450 569 -446
rect 657 -450 661 -446
rect 230 -462 234 -458
rect 284 -462 288 -458
rect 649 -460 653 -456
rect 332 -469 336 -465
rect 557 -466 561 -462
rect -75 -502 -71 -498
rect 49 -498 53 -494
rect 59 -491 63 -487
rect 565 -476 569 -472
rect 721 -479 725 -475
rect 731 -471 735 -467
rect 104 -505 108 -501
rect 241 -505 245 -501
rect 111 -515 115 -511
rect 669 -491 673 -487
rect 351 -507 355 -503
rect 234 -515 238 -511
rect -75 -538 -71 -534
rect 405 -512 409 -508
rect 481 -502 485 -498
rect 785 -481 789 -477
rect 854 -502 858 -498
rect 473 -512 477 -508
rect 546 -509 550 -505
rect 669 -509 673 -505
rect 326 -523 330 -519
rect 539 -519 543 -515
rect 676 -519 680 -515
rect 111 -533 115 -529
rect 496 -536 500 -532
rect 49 -553 53 -549
rect -6 -559 -2 -555
rect 59 -545 63 -541
rect 215 -548 219 -544
rect 721 -533 725 -529
rect 731 -526 735 -522
rect 854 -538 858 -534
rect 223 -558 227 -554
rect 131 -564 135 -560
rect 521 -552 525 -548
rect 123 -574 127 -570
rect 215 -574 219 -570
rect 405 -580 409 -576
rect 415 -587 419 -583
rect 785 -559 789 -555
rect 502 -590 506 -586
rect -106 -616 -102 -612
rect -96 -645 -92 -641
rect -80 -615 -76 -611
rect -70 -645 -66 -641
rect -50 -610 -46 -606
rect -20 -610 -16 -606
rect 104 -605 108 -601
rect 111 -615 115 -611
rect 200 -613 204 -609
rect 254 -613 258 -609
rect 364 -618 368 -614
rect 310 -624 314 -620
rect -40 -645 -36 -641
rect -10 -645 -6 -641
rect 111 -633 115 -629
rect 238 -632 242 -628
rect 184 -638 188 -634
rect 448 -606 452 -602
rect 458 -598 462 -594
rect 660 -592 664 -588
rect 474 -606 478 -602
rect 521 -606 525 -602
rect 294 -643 298 -639
rect 348 -643 352 -639
rect 572 -658 576 -654
rect 729 -613 733 -609
rect 799 -610 803 -606
rect 829 -610 833 -606
rect 789 -645 793 -641
rect 819 -645 823 -641
rect 859 -615 863 -611
rect 849 -645 853 -641
rect 885 -616 889 -612
rect 875 -645 879 -641
rect 224 -683 228 -679
rect 254 -683 258 -679
rect 190 -718 194 -714
rect 234 -718 238 -714
rect 264 -718 268 -714
rect 284 -683 288 -679
rect 294 -713 298 -709
rect 310 -683 314 -679
rect 464 -690 468 -686
rect 474 -698 478 -694
rect 591 -674 595 -670
rect 629 -670 633 -666
rect 320 -712 324 -708
rect 405 -717 409 -713
rect 415 -710 419 -706
rect 433 -710 437 -706
rect 220 -769 224 -765
rect 505 -717 509 -713
rect 515 -710 519 -706
rect 533 -710 537 -706
rect 639 -699 643 -695
rect 572 -712 576 -708
rect 655 -669 659 -665
rect 665 -699 669 -695
rect 685 -664 689 -660
rect 715 -664 719 -660
rect 759 -664 763 -660
rect 695 -699 699 -695
rect 725 -699 729 -695
rect 597 -728 601 -724
rect 390 -762 394 -758
rect 444 -762 448 -758
rect 397 -772 401 -768
rect 452 -772 456 -768
rect 289 -790 293 -786
rect 396 -825 400 -821
rect 310 -829 314 -825
rect 474 -825 478 -821
rect 345 -839 349 -835
rect 560 -829 564 -825
rect 525 -839 529 -835
rect 310 -859 314 -855
rect 560 -859 564 -855
rect 345 -869 349 -865
rect 525 -869 529 -865
rect 310 -889 314 -885
rect 417 -894 421 -890
rect 340 -899 344 -895
rect 453 -894 457 -890
rect 560 -889 564 -885
rect 530 -899 534 -895
rect 310 -915 314 -911
rect 560 -915 564 -911
rect 339 -925 343 -921
rect 531 -925 535 -921
<< metal1 >>
rect 278 -79 533 -76
rect 278 -94 282 -79
rect 271 -97 282 -94
rect 271 -106 274 -97
rect 278 -99 282 -97
rect 285 -92 293 -88
rect 307 -89 311 -82
rect 374 -85 437 -82
rect 374 -87 377 -85
rect 271 -109 282 -106
rect 278 -120 282 -109
rect 271 -123 282 -120
rect 271 -132 274 -123
rect 278 -125 282 -123
rect 285 -114 289 -92
rect 364 -92 371 -88
rect 384 -93 388 -85
rect 423 -93 427 -85
rect 434 -87 437 -85
rect 440 -92 447 -88
rect 500 -89 504 -82
rect 518 -92 526 -88
rect 303 -101 311 -97
rect 315 -101 324 -97
rect 487 -101 496 -97
rect 500 -101 508 -97
rect 308 -106 311 -101
rect 500 -106 503 -101
rect 308 -109 324 -106
rect 285 -118 293 -114
rect 308 -115 312 -109
rect 271 -135 282 -132
rect 278 -150 282 -135
rect 271 -153 282 -150
rect 271 -162 274 -153
rect 278 -155 282 -153
rect 285 -144 288 -118
rect 364 -118 371 -114
rect 392 -120 396 -113
rect 487 -109 503 -106
rect 415 -120 419 -113
rect 440 -118 447 -114
rect 499 -115 503 -109
rect 522 -114 526 -92
rect 529 -94 533 -79
rect 529 -97 540 -94
rect 529 -99 533 -97
rect 537 -106 540 -97
rect 518 -118 526 -114
rect 303 -127 307 -123
rect 364 -127 373 -123
rect 380 -124 385 -120
rect 378 -127 383 -124
rect 392 -125 397 -120
rect 414 -125 419 -120
rect 426 -124 431 -120
rect 304 -132 307 -127
rect 378 -132 381 -127
rect 428 -127 433 -124
rect 438 -127 447 -123
rect 504 -127 508 -123
rect 304 -135 324 -132
rect 364 -136 381 -132
rect 285 -148 292 -144
rect 313 -145 317 -143
rect 271 -165 282 -162
rect 278 -185 282 -165
rect 278 -195 282 -189
rect 285 -174 288 -148
rect 344 -147 356 -144
rect 344 -148 351 -147
rect 291 -157 292 -153
rect 324 -163 328 -156
rect 312 -166 328 -163
rect 363 -162 367 -153
rect 384 -159 388 -135
rect 423 -159 427 -135
rect 430 -132 433 -127
rect 504 -132 507 -127
rect 430 -136 447 -132
rect 487 -135 507 -132
rect 455 -147 467 -144
rect 460 -148 467 -147
rect 494 -145 498 -143
rect 523 -144 526 -118
rect 529 -109 540 -106
rect 529 -120 533 -109
rect 529 -123 540 -120
rect 529 -125 533 -123
rect 537 -132 540 -123
rect 519 -148 526 -144
rect 384 -162 427 -159
rect 285 -178 292 -174
rect 313 -175 317 -166
rect 285 -201 288 -178
rect 344 -178 351 -174
rect 291 -187 292 -183
rect 324 -193 328 -186
rect 371 -189 375 -182
rect 357 -193 364 -189
rect 312 -196 360 -193
rect 371 -194 376 -189
rect 285 -204 363 -201
rect 234 -207 288 -204
rect 363 -205 367 -204
rect 384 -205 388 -162
rect 234 -225 237 -207
rect 363 -208 388 -205
rect 252 -217 257 -216
rect 404 -217 407 -197
rect 423 -205 427 -162
rect 444 -162 448 -153
rect 483 -163 487 -156
rect 519 -157 520 -153
rect 483 -166 499 -163
rect 460 -178 467 -174
rect 494 -175 498 -166
rect 523 -174 526 -148
rect 529 -135 540 -132
rect 529 -150 533 -135
rect 529 -153 540 -150
rect 529 -155 533 -153
rect 537 -162 540 -153
rect 519 -178 526 -174
rect 436 -189 440 -182
rect 435 -194 440 -189
rect 447 -193 454 -189
rect 483 -193 487 -186
rect 519 -187 520 -183
rect 451 -196 499 -193
rect 523 -201 526 -178
rect 529 -165 540 -162
rect 529 -185 533 -165
rect 533 -189 572 -185
rect 448 -204 566 -201
rect 444 -205 448 -204
rect 423 -208 448 -205
rect 252 -221 264 -217
rect 333 -220 493 -217
rect 169 -229 242 -225
rect 333 -225 336 -220
rect 169 -246 172 -229
rect 253 -230 257 -228
rect 284 -229 336 -225
rect 250 -232 257 -230
rect 183 -238 188 -237
rect 241 -233 257 -232
rect 241 -235 253 -233
rect 183 -242 195 -238
rect 169 -250 173 -246
rect 155 -269 159 -262
rect 147 -296 151 -289
rect 141 -300 151 -296
rect 158 -300 164 -296
rect 147 -301 151 -300
rect 64 -308 69 -307
rect 57 -312 69 -308
rect 155 -312 159 -311
rect 173 -312 176 -250
rect 184 -253 188 -249
rect 215 -250 224 -246
rect 241 -249 245 -235
rect 292 -236 295 -229
rect 250 -249 254 -240
rect 290 -239 295 -236
rect 259 -249 263 -242
rect 285 -249 289 -242
rect 333 -247 336 -229
rect 370 -235 436 -232
rect 333 -251 343 -247
rect 370 -248 374 -235
rect 181 -256 188 -253
rect 181 -285 184 -256
rect 230 -262 233 -257
rect 199 -269 203 -262
rect 229 -269 233 -262
rect 333 -264 336 -251
rect 378 -241 415 -238
rect 363 -260 374 -256
rect 370 -265 374 -260
rect 378 -258 382 -241
rect 420 -241 429 -238
rect 403 -251 414 -247
rect 425 -248 429 -241
rect 407 -265 410 -251
rect 424 -260 429 -256
rect 425 -265 429 -260
rect 432 -258 436 -235
rect 490 -247 493 -220
rect 563 -225 566 -204
rect 569 -218 572 -189
rect 581 -214 596 -211
rect 581 -218 584 -214
rect 593 -218 596 -214
rect 607 -214 622 -211
rect 607 -218 610 -214
rect 619 -218 622 -214
rect 637 -214 652 -211
rect 637 -218 640 -214
rect 649 -218 652 -214
rect 569 -222 586 -218
rect 593 -222 612 -218
rect 619 -222 642 -218
rect 649 -222 672 -218
rect 676 -222 684 -218
rect 563 -228 691 -225
rect 575 -229 605 -228
rect 575 -233 579 -229
rect 601 -233 605 -229
rect 631 -232 635 -228
rect 640 -232 644 -231
rect 661 -232 665 -228
rect 670 -232 674 -231
rect 688 -238 691 -228
rect 483 -251 511 -247
rect 573 -251 576 -247
rect 584 -248 588 -243
rect 610 -244 614 -243
rect 688 -241 709 -238
rect 610 -247 622 -244
rect 584 -251 602 -248
rect 593 -252 602 -251
rect 584 -264 588 -255
rect 336 -269 343 -265
rect 370 -269 383 -265
rect 407 -266 414 -265
rect 370 -276 374 -269
rect 411 -269 414 -266
rect 425 -269 443 -265
rect 593 -264 596 -252
rect 619 -264 622 -247
rect 650 -253 653 -252
rect 630 -257 632 -253
rect 650 -257 662 -253
rect 650 -264 653 -257
rect 680 -264 683 -252
rect 643 -268 653 -264
rect 673 -268 683 -264
rect 425 -275 429 -269
rect 302 -279 374 -276
rect 181 -289 191 -285
rect 211 -289 221 -285
rect 181 -301 184 -289
rect 211 -296 214 -289
rect 202 -300 214 -296
rect 232 -300 234 -296
rect 211 -301 214 -300
rect 242 -306 245 -289
rect 268 -301 271 -289
rect 276 -298 280 -289
rect 262 -302 271 -301
rect 262 -305 280 -302
rect 242 -309 254 -306
rect 155 -315 176 -312
rect 250 -310 254 -309
rect 276 -310 280 -305
rect 288 -306 290 -302
rect 26 -320 37 -316
rect 155 -316 159 -315
rect 26 -327 29 -320
rect 64 -321 68 -319
rect 79 -320 159 -316
rect 64 -323 71 -321
rect 64 -324 80 -323
rect 68 -326 80 -324
rect 26 -330 31 -327
rect 32 -340 36 -333
rect 58 -340 62 -333
rect 67 -340 71 -331
rect 76 -340 80 -326
rect 133 -329 138 -328
rect 126 -333 138 -329
rect 97 -341 106 -337
rect 149 -337 152 -320
rect 173 -325 176 -315
rect 190 -322 194 -321
rect 199 -325 203 -321
rect 220 -322 224 -321
rect 229 -325 233 -321
rect 259 -324 263 -320
rect 285 -324 289 -320
rect 259 -325 289 -324
rect 173 -328 289 -325
rect 133 -344 137 -340
rect 148 -341 152 -337
rect 180 -334 188 -331
rect 133 -347 140 -344
rect 88 -353 91 -348
rect 88 -360 92 -353
rect 118 -360 122 -353
rect 137 -376 140 -347
rect -101 -387 -86 -384
rect -101 -391 -98 -387
rect -89 -391 -86 -387
rect -75 -387 -60 -384
rect -75 -391 -72 -387
rect -63 -391 -60 -387
rect -45 -387 -30 -384
rect -45 -391 -42 -387
rect -33 -391 -30 -387
rect 41 -389 45 -380
rect 100 -380 110 -376
rect 130 -380 140 -376
rect -119 -395 -96 -391
rect -89 -395 -70 -391
rect -63 -395 -40 -391
rect -33 -395 -10 -391
rect -6 -395 15 -391
rect 50 -392 53 -380
rect -119 -641 -116 -395
rect -107 -401 9 -398
rect -107 -402 -77 -401
rect -107 -406 -103 -402
rect -81 -406 -77 -402
rect -51 -405 -47 -401
rect -42 -405 -38 -404
rect -21 -405 -17 -401
rect -12 -405 -8 -404
rect -113 -424 -106 -420
rect -98 -421 -94 -416
rect -72 -417 -68 -416
rect -72 -420 -60 -417
rect -98 -424 -80 -421
rect -89 -425 -80 -424
rect -98 -437 -94 -428
rect -89 -437 -86 -425
rect -63 -437 -60 -420
rect -32 -426 -29 -425
rect -52 -430 -50 -426
rect -32 -430 -20 -426
rect -32 -437 -29 -430
rect -2 -437 1 -425
rect -39 -441 -29 -437
rect -9 -441 1 -437
rect -51 -464 -47 -457
rect -21 -464 -17 -457
rect -51 -469 -48 -464
rect -2 -470 1 -441
rect -6 -473 1 -470
rect -107 -484 -103 -477
rect -81 -484 -77 -477
rect -113 -490 -108 -487
rect -72 -486 -68 -477
rect -113 -497 -110 -490
rect -63 -491 -59 -477
rect -42 -480 -33 -476
rect -6 -477 -2 -473
rect 6 -476 9 -401
rect 12 -430 15 -395
rect 50 -393 59 -392
rect 30 -397 33 -393
rect 41 -396 59 -393
rect 41 -401 45 -396
rect 76 -397 79 -380
rect 107 -387 110 -380
rect 87 -391 89 -387
rect 107 -391 119 -387
rect 107 -392 110 -391
rect 137 -392 140 -380
rect 67 -400 79 -397
rect 67 -401 71 -400
rect 32 -415 36 -411
rect 58 -415 62 -411
rect 32 -416 62 -415
rect 88 -416 92 -412
rect 97 -413 101 -412
rect 118 -416 122 -412
rect 127 -413 131 -412
rect 145 -416 148 -341
rect 32 -419 148 -416
rect 38 -426 43 -422
rect 64 -426 69 -422
rect 94 -426 99 -422
rect 124 -426 129 -422
rect 38 -430 41 -426
rect 64 -430 67 -426
rect 94 -430 97 -426
rect 124 -430 127 -426
rect 180 -430 183 -334
rect 192 -335 215 -331
rect 222 -335 245 -331
rect 252 -335 271 -331
rect 278 -335 283 -331
rect 212 -339 215 -335
rect 224 -339 227 -335
rect 212 -342 227 -339
rect 242 -339 245 -335
rect 254 -339 257 -335
rect 242 -342 257 -339
rect 268 -339 271 -335
rect 280 -338 283 -335
rect 268 -342 278 -339
rect 302 -346 305 -279
rect 325 -283 359 -282
rect 328 -285 359 -283
rect 337 -292 341 -285
rect 355 -292 359 -285
rect 346 -319 350 -312
rect 367 -319 370 -279
rect 489 -279 506 -276
rect 386 -284 418 -281
rect 386 -311 390 -284
rect 414 -291 418 -284
rect 432 -285 482 -282
rect 432 -291 435 -285
rect 418 -295 435 -291
rect 223 -349 305 -346
rect 308 -322 350 -319
rect 223 -376 226 -349
rect 308 -355 311 -322
rect 284 -358 311 -355
rect 284 -367 288 -358
rect 277 -371 289 -367
rect 300 -368 304 -366
rect 12 -433 183 -430
rect 186 -379 226 -376
rect 20 -476 23 -468
rect 186 -475 189 -379
rect 246 -380 250 -378
rect 277 -379 289 -375
rect 284 -380 289 -379
rect 300 -380 304 -372
rect 284 -386 289 -385
rect 222 -390 235 -386
rect 277 -390 289 -386
rect 9 -480 13 -476
rect -13 -488 -1 -484
rect -71 -493 -59 -491
rect -75 -494 -59 -493
rect -6 -489 -1 -488
rect -75 -496 -68 -494
rect -113 -501 -102 -497
rect -75 -498 -71 -496
rect 10 -497 13 -480
rect -113 -535 -110 -501
rect -60 -501 13 -497
rect -82 -509 -70 -505
rect -75 -510 -70 -509
rect 10 -512 13 -501
rect 20 -480 48 -476
rect -75 -527 -70 -526
rect -82 -531 -70 -527
rect -113 -539 -102 -535
rect 10 -535 13 -517
rect -113 -546 -110 -539
rect -75 -540 -71 -538
rect -60 -539 13 -535
rect -75 -542 -68 -540
rect -75 -543 -59 -542
rect -71 -545 -59 -543
rect -113 -549 -108 -546
rect -107 -559 -103 -552
rect -81 -559 -77 -552
rect -72 -559 -68 -550
rect -63 -559 -59 -545
rect -6 -548 -1 -547
rect -13 -552 -1 -548
rect -42 -560 -33 -556
rect 10 -556 13 -539
rect -6 -563 -2 -559
rect 9 -560 13 -556
rect -6 -566 1 -563
rect -51 -572 -48 -567
rect -51 -579 -47 -572
rect -21 -579 -17 -572
rect -2 -595 1 -566
rect -98 -608 -94 -599
rect -39 -599 -29 -595
rect -9 -599 1 -595
rect -89 -611 -86 -599
rect -89 -612 -80 -611
rect -113 -616 -106 -612
rect -98 -615 -80 -612
rect -98 -620 -94 -615
rect -63 -616 -60 -599
rect -32 -606 -29 -599
rect -52 -610 -50 -606
rect -32 -610 -20 -606
rect -32 -611 -29 -610
rect -2 -611 1 -599
rect -72 -619 -60 -616
rect -72 -620 -68 -619
rect -107 -634 -103 -630
rect -81 -634 -77 -630
rect -107 -635 -77 -634
rect -51 -635 -47 -631
rect -42 -632 -38 -631
rect -21 -635 -17 -631
rect -12 -632 -8 -631
rect 6 -635 9 -560
rect 20 -587 23 -480
rect 33 -491 59 -487
rect 33 -549 36 -491
rect 66 -494 70 -480
rect 111 -478 189 -475
rect 192 -398 202 -394
rect 192 -459 195 -398
rect 230 -405 234 -397
rect 241 -413 245 -398
rect 257 -405 261 -398
rect 284 -402 288 -397
rect 299 -398 300 -394
rect 308 -402 311 -358
rect 331 -360 334 -322
rect 337 -332 341 -322
rect 358 -323 370 -319
rect 479 -321 482 -285
rect 348 -331 368 -327
rect 365 -338 368 -331
rect 378 -338 382 -331
rect 396 -338 400 -331
rect 479 -333 483 -326
rect 365 -342 382 -338
rect 389 -342 400 -338
rect 407 -342 425 -338
rect 378 -343 382 -342
rect 396 -345 400 -342
rect 396 -349 409 -345
rect 417 -349 426 -345
rect 355 -354 359 -352
rect 355 -357 372 -354
rect 386 -354 390 -353
rect 405 -350 409 -349
rect 377 -357 390 -354
rect 331 -363 383 -360
rect 380 -370 383 -363
rect 386 -364 390 -357
rect 396 -364 400 -360
rect 414 -364 418 -360
rect 386 -367 418 -364
rect 284 -405 311 -402
rect 241 -416 317 -413
rect 284 -423 311 -420
rect 284 -432 288 -423
rect 277 -436 289 -432
rect 300 -433 304 -431
rect 246 -445 250 -443
rect 277 -444 289 -440
rect 284 -445 289 -444
rect 300 -445 304 -437
rect 284 -451 289 -450
rect 222 -455 235 -451
rect 277 -455 289 -451
rect 192 -463 202 -459
rect 39 -498 49 -494
rect 57 -498 78 -494
rect 83 -497 108 -494
rect 39 -503 42 -498
rect 57 -499 61 -498
rect 86 -504 93 -500
rect 104 -501 108 -497
rect 39 -541 42 -508
rect 48 -512 52 -509
rect 66 -513 70 -509
rect 86 -513 89 -504
rect 103 -513 108 -509
rect 53 -516 89 -513
rect 48 -520 52 -517
rect 86 -518 89 -516
rect 104 -518 108 -513
rect 111 -511 114 -478
rect 192 -486 195 -463
rect 230 -470 234 -462
rect 241 -481 245 -463
rect 257 -470 261 -463
rect 284 -466 288 -462
rect 299 -463 300 -459
rect 308 -467 311 -423
rect 289 -470 311 -467
rect 314 -481 317 -416
rect 352 -421 356 -414
rect 344 -454 348 -441
rect 355 -453 363 -449
rect 387 -453 390 -367
rect 372 -456 390 -453
rect 372 -458 375 -456
rect 356 -463 370 -460
rect 356 -464 375 -463
rect 336 -469 338 -465
rect 356 -480 363 -476
rect 241 -484 317 -481
rect 169 -489 195 -486
rect 169 -500 172 -489
rect 162 -504 187 -500
rect 86 -522 93 -518
rect 104 -522 122 -518
rect 86 -528 89 -522
rect 86 -532 93 -528
rect 98 -532 100 -528
rect 111 -529 115 -522
rect 169 -528 172 -504
rect 142 -532 172 -528
rect 110 -540 122 -536
rect 39 -545 59 -541
rect 66 -549 70 -540
rect 111 -547 115 -540
rect 178 -543 181 -504
rect 234 -511 238 -494
rect 242 -497 243 -494
rect 241 -501 245 -497
rect 257 -500 260 -484
rect 256 -504 263 -500
rect 325 -503 329 -496
rect 241 -513 246 -509
rect 241 -518 245 -513
rect 260 -518 263 -504
rect 313 -507 329 -503
rect 227 -522 245 -518
rect 256 -522 259 -518
rect 241 -527 245 -522
rect 215 -532 240 -529
rect 313 -527 316 -507
rect 325 -508 329 -507
rect 333 -503 337 -496
rect 344 -503 348 -496
rect 333 -508 338 -503
rect 343 -508 348 -503
rect 355 -507 363 -503
rect 360 -508 363 -507
rect 393 -508 396 -386
rect 423 -446 426 -349
rect 471 -366 475 -353
rect 482 -365 490 -361
rect 503 -372 506 -279
rect 631 -291 635 -284
rect 661 -291 665 -284
rect 631 -296 634 -291
rect 680 -297 683 -268
rect 676 -300 683 -297
rect 575 -311 579 -304
rect 601 -311 605 -304
rect 569 -317 574 -314
rect 610 -313 614 -304
rect 569 -321 572 -317
rect 619 -318 623 -304
rect 640 -307 649 -303
rect 676 -304 680 -300
rect 688 -303 691 -241
rect 705 -242 709 -241
rect 713 -253 717 -252
rect 700 -257 706 -253
rect 713 -257 723 -253
rect 713 -264 717 -257
rect 781 -261 786 -260
rect 774 -265 786 -261
rect 743 -273 754 -269
rect 743 -280 746 -273
rect 781 -274 785 -272
rect 796 -273 864 -269
rect 781 -276 788 -274
rect 781 -277 797 -276
rect 785 -279 797 -277
rect 743 -283 748 -280
rect 705 -291 709 -284
rect 724 -286 748 -283
rect 724 -291 727 -286
rect 709 -294 727 -291
rect 749 -293 753 -286
rect 775 -293 779 -286
rect 784 -293 788 -284
rect 793 -293 797 -279
rect 850 -282 855 -281
rect 843 -286 855 -282
rect 814 -294 823 -290
rect 866 -290 869 -274
rect 850 -297 854 -293
rect 865 -294 869 -290
rect 850 -300 857 -297
rect 691 -307 695 -303
rect 669 -315 681 -311
rect 611 -320 623 -318
rect 518 -324 572 -321
rect 607 -321 623 -320
rect 676 -316 681 -315
rect 607 -323 614 -321
rect 692 -323 695 -307
rect 805 -306 808 -301
rect 805 -313 809 -306
rect 835 -313 839 -306
rect 569 -328 580 -324
rect 607 -325 611 -323
rect 622 -328 690 -324
rect 854 -329 857 -300
rect 600 -336 612 -332
rect 607 -337 612 -336
rect 758 -342 762 -333
rect 817 -333 827 -329
rect 847 -333 857 -329
rect 767 -345 770 -333
rect 767 -346 776 -345
rect 649 -350 750 -346
rect 758 -349 776 -346
rect 649 -354 653 -350
rect 758 -354 762 -349
rect 793 -350 796 -333
rect 824 -340 827 -333
rect 804 -344 806 -340
rect 824 -344 836 -340
rect 824 -345 827 -344
rect 854 -345 857 -333
rect 612 -358 622 -354
rect 649 -358 662 -354
rect 784 -353 796 -350
rect 784 -354 788 -353
rect 862 -356 865 -294
rect 879 -313 883 -306
rect 887 -340 891 -333
rect 874 -344 880 -340
rect 887 -344 897 -340
rect 887 -345 891 -344
rect 879 -356 883 -355
rect 612 -360 615 -358
rect 649 -363 653 -358
rect 862 -359 883 -356
rect 545 -369 606 -366
rect 483 -376 523 -372
rect 545 -376 549 -369
rect 463 -381 465 -377
rect 520 -384 523 -376
rect 544 -380 556 -376
rect 603 -378 606 -369
rect 612 -372 615 -365
rect 642 -367 653 -363
rect 612 -375 622 -372
rect 603 -381 612 -378
rect 609 -383 612 -381
rect 649 -383 653 -375
rect 520 -388 534 -384
rect 483 -392 490 -388
rect 520 -394 523 -388
rect 545 -394 549 -387
rect 576 -388 606 -384
rect 609 -386 653 -383
rect 520 -398 527 -394
rect 538 -398 556 -394
rect 452 -415 456 -408
rect 440 -419 456 -415
rect 440 -439 443 -419
rect 452 -420 456 -419
rect 460 -415 464 -408
rect 471 -415 475 -408
rect 520 -412 523 -398
rect 538 -403 542 -398
rect 537 -407 542 -403
rect 460 -420 465 -415
rect 470 -420 475 -415
rect 482 -419 487 -415
rect 523 -416 527 -412
rect 479 -431 483 -430
rect 451 -435 453 -431
rect 457 -435 465 -431
rect 487 -439 490 -420
rect 440 -442 490 -439
rect 538 -441 542 -415
rect 545 -423 549 -405
rect 603 -412 606 -388
rect 657 -387 661 -365
rect 749 -368 753 -364
rect 775 -368 779 -364
rect 749 -369 779 -368
rect 805 -369 809 -365
rect 814 -366 818 -365
rect 835 -369 839 -365
rect 844 -366 848 -365
rect 862 -367 865 -359
rect 749 -371 860 -369
rect 750 -372 860 -371
rect 682 -376 690 -372
rect 657 -390 673 -387
rect 669 -398 673 -390
rect 692 -398 695 -378
rect 747 -379 760 -375
rect 767 -379 786 -375
rect 793 -379 816 -375
rect 824 -379 846 -375
rect 755 -383 758 -379
rect 767 -383 770 -379
rect 755 -386 770 -383
rect 781 -383 784 -379
rect 793 -383 796 -379
rect 781 -386 796 -383
rect 812 -383 815 -379
rect 824 -383 828 -379
rect 812 -387 828 -383
rect 812 -391 815 -387
rect 824 -391 828 -387
rect 843 -387 858 -384
rect 843 -391 846 -387
rect 855 -391 858 -387
rect 869 -387 884 -384
rect 869 -391 872 -387
rect 881 -391 884 -387
rect 793 -395 815 -391
rect 823 -395 846 -391
rect 853 -395 872 -391
rect 879 -395 902 -391
rect 662 -402 680 -398
rect 691 -402 698 -398
rect 596 -416 603 -412
rect 608 -416 615 -414
rect 608 -417 622 -416
rect 612 -420 622 -417
rect 669 -427 673 -409
rect 676 -407 680 -402
rect 676 -411 681 -407
rect 565 -430 673 -427
rect 695 -416 698 -402
rect 565 -439 569 -430
rect 676 -433 680 -419
rect 691 -420 698 -416
rect 774 -401 860 -398
rect 654 -436 680 -433
rect 649 -439 654 -438
rect 523 -444 542 -441
rect 564 -443 576 -439
rect 612 -443 622 -439
rect 649 -443 662 -439
rect 523 -446 526 -444
rect 423 -449 526 -446
rect 404 -481 408 -461
rect 412 -508 416 -501
rect 423 -508 426 -449
rect 529 -451 554 -447
rect 439 -471 442 -457
rect 360 -511 405 -508
rect 352 -519 356 -518
rect 324 -523 326 -519
rect 330 -523 338 -519
rect 360 -527 363 -511
rect 313 -530 363 -527
rect 393 -512 405 -511
rect 412 -512 426 -508
rect 429 -474 442 -471
rect 178 -547 188 -543
rect 215 -544 219 -532
rect 393 -535 396 -512
rect 412 -513 416 -512
rect 33 -553 49 -549
rect 57 -553 77 -549
rect 57 -560 61 -553
rect 111 -550 135 -547
rect 82 -553 108 -550
rect 105 -556 127 -553
rect 89 -563 93 -559
rect 98 -563 102 -559
rect 48 -587 52 -580
rect 66 -587 70 -580
rect 20 -590 65 -587
rect 89 -600 92 -563
rect 123 -570 127 -556
rect 131 -560 135 -550
rect 162 -563 172 -559
rect 169 -566 172 -563
rect 178 -561 181 -547
rect 223 -538 396 -535
rect 208 -556 219 -552
rect 215 -561 219 -556
rect 223 -554 227 -538
rect 248 -547 252 -543
rect 178 -565 188 -561
rect 215 -565 228 -561
rect 178 -566 181 -565
rect 131 -572 142 -568
rect 181 -571 188 -569
rect 131 -577 135 -572
rect 169 -577 172 -571
rect 178 -573 188 -571
rect 215 -570 219 -565
rect 252 -569 255 -547
rect 272 -547 390 -544
rect 404 -558 408 -523
rect 429 -550 432 -474
rect 436 -491 439 -484
rect 473 -491 477 -460
rect 529 -472 532 -451
rect 565 -455 569 -450
rect 596 -451 603 -447
rect 603 -455 606 -451
rect 556 -459 569 -455
rect 596 -458 606 -455
rect 612 -457 615 -443
rect 649 -448 653 -443
rect 642 -452 653 -448
rect 612 -458 622 -457
rect 596 -459 622 -458
rect 533 -477 536 -473
rect 557 -482 561 -466
rect 565 -464 569 -459
rect 603 -461 622 -459
rect 565 -468 576 -464
rect 526 -485 561 -482
rect 603 -473 606 -466
rect 565 -488 569 -476
rect 596 -477 606 -473
rect 539 -491 569 -488
rect 612 -488 615 -461
rect 649 -470 653 -460
rect 657 -464 661 -450
rect 692 -457 695 -420
rect 718 -433 763 -430
rect 714 -440 718 -433
rect 732 -440 736 -433
rect 682 -461 683 -457
rect 688 -460 695 -457
rect 657 -467 679 -464
rect 676 -470 702 -467
rect 649 -473 673 -470
rect 723 -467 727 -460
rect 707 -471 727 -467
rect 735 -471 751 -467
rect 669 -480 673 -473
rect 714 -480 718 -471
rect 725 -479 745 -475
rect 662 -484 674 -480
rect 436 -495 446 -491
rect 473 -495 486 -491
rect 436 -509 439 -495
rect 473 -500 477 -495
rect 539 -498 544 -496
rect 612 -492 642 -488
rect 466 -504 477 -500
rect 436 -513 446 -509
rect 473 -542 477 -512
rect 481 -516 485 -502
rect 523 -502 528 -498
rect 539 -502 557 -498
rect 523 -503 524 -502
rect 521 -509 524 -503
rect 539 -507 543 -502
rect 506 -513 524 -509
rect 538 -511 543 -507
rect 521 -516 524 -513
rect 521 -520 528 -516
rect 483 -528 533 -525
rect 483 -548 486 -528
rect 494 -536 496 -532
rect 500 -536 508 -532
rect 530 -533 533 -528
rect 522 -537 526 -536
rect 530 -538 531 -533
rect 539 -534 542 -519
rect 546 -525 550 -509
rect 612 -516 615 -492
rect 669 -498 673 -491
rect 684 -492 698 -488
rect 695 -498 698 -492
rect 662 -502 680 -498
rect 691 -502 698 -498
rect 597 -520 622 -516
rect 539 -537 548 -534
rect 495 -548 499 -547
rect 429 -553 442 -550
rect 483 -552 499 -548
rect 230 -573 255 -569
rect 122 -580 135 -577
rect 122 -581 127 -580
rect 104 -585 127 -584
rect 132 -585 135 -580
rect 162 -581 172 -577
rect 208 -581 220 -577
rect 104 -587 135 -585
rect -107 -638 9 -635
rect 86 -604 93 -600
rect 104 -601 108 -587
rect 215 -590 219 -581
rect 252 -586 255 -573
rect 378 -561 384 -558
rect 378 -586 381 -561
rect 389 -561 422 -558
rect 404 -565 408 -561
rect 422 -565 426 -561
rect 413 -576 417 -575
rect 86 -618 89 -604
rect 111 -593 219 -590
rect 243 -589 381 -586
rect 386 -579 405 -576
rect 386 -587 389 -579
rect 401 -580 405 -579
rect 413 -580 436 -576
rect 398 -587 415 -583
rect 103 -613 108 -609
rect 104 -618 108 -613
rect 111 -611 115 -593
rect 162 -604 169 -600
rect 177 -604 204 -601
rect 86 -622 93 -618
rect 104 -622 122 -618
rect 86 -628 89 -622
rect 86 -632 100 -628
rect 111 -629 115 -622
rect 169 -627 172 -604
rect -119 -645 -96 -641
rect -89 -645 -70 -641
rect -63 -645 -40 -641
rect -33 -645 -10 -641
rect -101 -649 -98 -645
rect -89 -649 -86 -645
rect -101 -652 -86 -649
rect -75 -649 -72 -645
rect -63 -649 -60 -645
rect -75 -652 -60 -649
rect -45 -649 -42 -645
rect -33 -649 -30 -645
rect -45 -652 -30 -649
rect 86 -659 89 -632
rect 142 -632 169 -628
rect 110 -640 122 -636
rect 111 -643 115 -640
rect 177 -646 180 -604
rect 188 -612 189 -608
rect 200 -609 204 -604
rect 227 -608 231 -601
rect 243 -608 247 -589
rect 254 -609 258 -601
rect 293 -605 304 -602
rect 348 -604 375 -601
rect 293 -608 296 -605
rect 286 -612 296 -608
rect 199 -620 211 -616
rect 253 -620 266 -616
rect 199 -621 204 -620
rect 184 -634 188 -626
rect 199 -627 204 -626
rect 291 -621 294 -612
rect 348 -613 352 -604
rect 341 -617 353 -613
rect 364 -614 368 -612
rect 273 -624 294 -621
rect 199 -631 211 -627
rect 238 -628 242 -626
rect 273 -628 276 -624
rect 310 -626 314 -624
rect 341 -625 353 -621
rect 256 -631 276 -628
rect 184 -640 188 -638
rect 199 -639 211 -635
rect 200 -648 204 -639
rect 180 -651 204 -648
rect 256 -640 259 -631
rect 348 -626 353 -625
rect 364 -626 368 -618
rect 348 -632 353 -631
rect 286 -636 299 -632
rect 341 -636 353 -632
rect 256 -644 266 -640
rect 256 -651 259 -644
rect 294 -651 298 -643
rect 86 -662 208 -659
rect 305 -659 309 -644
rect 321 -651 325 -644
rect 348 -648 352 -643
rect 363 -644 364 -640
rect 372 -648 375 -604
rect 348 -651 370 -648
rect 378 -659 381 -589
rect 422 -594 426 -580
rect 433 -602 436 -580
rect 439 -594 442 -553
rect 495 -559 499 -552
rect 503 -552 508 -547
rect 513 -552 518 -547
rect 530 -548 533 -538
rect 525 -552 533 -548
rect 503 -559 507 -552
rect 514 -559 518 -552
rect 447 -569 468 -566
rect 447 -573 451 -569
rect 439 -598 458 -594
rect 465 -602 469 -593
rect 473 -591 477 -566
rect 526 -579 533 -575
rect 506 -590 508 -586
rect 526 -595 542 -591
rect 481 -602 485 -601
rect 433 -606 448 -602
rect 456 -606 474 -602
rect 481 -606 497 -602
rect 456 -613 460 -606
rect 481 -613 485 -606
rect 404 -643 408 -634
rect 447 -640 451 -633
rect 465 -640 469 -633
rect 473 -640 477 -633
rect 447 -643 472 -640
rect 213 -662 381 -659
rect 404 -649 408 -648
rect 463 -649 466 -643
rect 404 -652 481 -649
rect 404 -659 408 -652
rect 83 -668 393 -665
rect 248 -675 263 -672
rect 248 -679 251 -675
rect 260 -679 263 -675
rect 278 -675 293 -672
rect 278 -679 281 -675
rect 290 -679 293 -675
rect 304 -675 319 -672
rect 304 -679 307 -675
rect 316 -679 319 -675
rect 228 -683 251 -679
rect 258 -683 281 -679
rect 288 -683 307 -679
rect 314 -683 338 -679
rect 213 -689 325 -686
rect 209 -699 212 -690
rect 226 -693 230 -692
rect 235 -693 239 -689
rect 256 -693 260 -692
rect 265 -693 269 -689
rect 295 -690 325 -689
rect 295 -694 299 -690
rect 321 -694 325 -690
rect 191 -702 212 -699
rect 191 -703 195 -702
rect 183 -714 187 -713
rect 177 -718 187 -714
rect 194 -718 200 -714
rect 183 -725 187 -718
rect 191 -752 195 -745
rect 209 -764 212 -702
rect 286 -705 290 -704
rect 278 -708 290 -705
rect 217 -725 220 -713
rect 247 -714 250 -713
rect 238 -718 250 -714
rect 268 -718 270 -714
rect 247 -725 250 -718
rect 278 -725 281 -708
rect 312 -709 316 -704
rect 298 -712 316 -709
rect 324 -712 327 -708
rect 298 -713 307 -712
rect 304 -725 307 -713
rect 217 -729 227 -725
rect 247 -729 257 -725
rect 312 -725 316 -716
rect 335 -718 338 -683
rect 390 -707 393 -668
rect 432 -679 436 -652
rect 463 -659 467 -652
rect 481 -659 485 -652
rect 472 -686 476 -679
rect 451 -690 464 -686
rect 472 -690 491 -686
rect 422 -706 426 -699
rect 440 -706 444 -699
rect 451 -706 454 -690
rect 390 -710 415 -707
rect 422 -710 433 -706
rect 440 -710 454 -706
rect 457 -698 474 -694
rect 422 -713 426 -710
rect 333 -721 338 -718
rect 398 -717 405 -713
rect 413 -717 426 -713
rect 440 -711 444 -710
rect 457 -713 460 -698
rect 481 -699 485 -690
rect 454 -716 460 -713
rect 488 -713 491 -690
rect 494 -706 497 -606
rect 514 -614 518 -601
rect 525 -606 531 -602
rect 539 -628 542 -595
rect 522 -641 526 -634
rect 545 -637 548 -537
rect 571 -600 575 -520
rect 670 -531 673 -509
rect 676 -507 680 -502
rect 695 -504 698 -502
rect 732 -503 736 -500
rect 676 -511 681 -507
rect 695 -508 709 -504
rect 714 -507 731 -504
rect 695 -516 698 -508
rect 714 -511 718 -507
rect 732 -511 736 -508
rect 742 -512 745 -479
rect 676 -523 680 -519
rect 691 -520 698 -516
rect 723 -522 727 -521
rect 742 -522 745 -517
rect 676 -526 701 -523
rect 706 -526 727 -522
rect 735 -526 745 -522
rect 748 -485 751 -471
rect 748 -490 752 -485
rect 617 -534 673 -531
rect 571 -616 575 -605
rect 552 -619 575 -616
rect 522 -649 526 -646
rect 552 -649 555 -619
rect 571 -626 575 -619
rect 504 -652 555 -649
rect 504 -659 508 -652
rect 532 -679 536 -652
rect 565 -658 572 -654
rect 579 -659 583 -646
rect 557 -669 571 -665
rect 589 -674 591 -670
rect 564 -685 571 -681
rect 522 -706 526 -699
rect 540 -706 544 -699
rect 494 -710 515 -706
rect 522 -710 533 -706
rect 540 -709 561 -706
rect 579 -708 583 -701
rect 590 -708 594 -701
rect 540 -710 572 -709
rect 522 -713 526 -710
rect 217 -758 220 -729
rect 235 -752 239 -745
rect 265 -752 269 -745
rect 266 -757 269 -752
rect 217 -761 224 -758
rect 205 -768 209 -764
rect 220 -765 224 -761
rect 205 -785 208 -768
rect 251 -768 260 -764
rect 219 -776 231 -772
rect 219 -777 224 -776
rect 277 -779 281 -765
rect 286 -774 290 -765
rect 295 -772 299 -765
rect 321 -772 325 -765
rect 326 -778 330 -775
rect 277 -781 289 -779
rect 277 -782 293 -781
rect 286 -784 293 -782
rect 205 -789 278 -785
rect 289 -786 293 -784
rect 327 -785 330 -778
rect 320 -789 330 -785
rect 288 -797 300 -793
rect 288 -798 293 -797
rect 333 -804 336 -721
rect 398 -738 401 -717
rect 413 -718 417 -717
rect 404 -732 408 -728
rect 422 -732 426 -728
rect 432 -730 436 -721
rect 404 -735 431 -732
rect 397 -751 401 -743
rect 416 -751 419 -735
rect 454 -736 457 -716
rect 488 -717 505 -713
rect 513 -717 526 -713
rect 540 -711 544 -710
rect 558 -712 572 -710
rect 463 -730 467 -719
rect 513 -718 517 -717
rect 504 -732 508 -728
rect 522 -732 526 -728
rect 532 -732 536 -721
rect 467 -735 552 -732
rect 564 -732 567 -712
rect 579 -713 584 -708
rect 589 -713 594 -708
rect 598 -708 602 -701
rect 598 -712 614 -708
rect 598 -713 602 -712
rect 571 -724 575 -723
rect 589 -728 597 -724
rect 601 -728 603 -724
rect 611 -732 614 -712
rect 564 -735 614 -732
rect 453 -738 457 -736
rect 617 -738 620 -534
rect 714 -540 718 -526
rect 748 -529 751 -490
rect 725 -533 751 -529
rect 760 -540 763 -433
rect 774 -476 777 -401
rect 791 -405 795 -404
rect 800 -405 804 -401
rect 821 -405 825 -404
rect 830 -405 834 -401
rect 866 -402 890 -398
rect 860 -406 864 -404
rect 886 -406 890 -402
rect 851 -417 855 -416
rect 843 -420 855 -417
rect 782 -437 785 -425
rect 812 -426 815 -425
rect 803 -430 815 -426
rect 833 -430 835 -426
rect 812 -437 815 -430
rect 843 -437 846 -420
rect 877 -421 881 -416
rect 863 -424 881 -421
rect 889 -424 896 -420
rect 863 -425 872 -424
rect 869 -437 872 -425
rect 782 -441 792 -437
rect 812 -441 822 -437
rect 877 -437 881 -428
rect 782 -470 785 -441
rect 800 -464 804 -457
rect 830 -464 834 -457
rect 831 -469 834 -464
rect 782 -473 789 -470
rect 770 -480 774 -476
rect 785 -477 789 -473
rect 770 -497 773 -480
rect 816 -480 825 -476
rect 784 -488 796 -484
rect 784 -489 789 -488
rect 842 -491 846 -477
rect 851 -486 855 -477
rect 860 -484 864 -477
rect 886 -484 890 -477
rect 891 -490 896 -487
rect 842 -493 854 -491
rect 842 -494 858 -493
rect 851 -496 858 -494
rect 770 -498 843 -497
rect 775 -501 843 -498
rect 854 -498 858 -496
rect 893 -497 896 -490
rect 885 -501 896 -497
rect 736 -544 763 -540
rect 760 -568 763 -544
rect 770 -535 773 -503
rect 853 -509 865 -505
rect 853 -510 858 -509
rect 853 -527 858 -526
rect 853 -531 865 -527
rect 770 -539 843 -535
rect 893 -535 896 -501
rect 770 -556 773 -539
rect 854 -540 858 -538
rect 885 -539 896 -535
rect 851 -542 858 -540
rect 784 -548 789 -547
rect 842 -543 858 -542
rect 842 -545 854 -543
rect 784 -552 796 -548
rect 770 -560 774 -556
rect 660 -581 665 -580
rect 653 -585 665 -581
rect 623 -593 633 -589
rect 774 -589 777 -560
rect 785 -563 789 -559
rect 816 -560 825 -556
rect 842 -559 846 -545
rect 893 -546 896 -539
rect 851 -559 855 -550
rect 891 -549 896 -546
rect 860 -559 864 -552
rect 886 -559 890 -552
rect 623 -600 626 -593
rect 660 -594 664 -592
rect 675 -593 777 -589
rect 660 -596 667 -594
rect 660 -597 676 -596
rect 664 -599 676 -597
rect 623 -603 627 -600
rect 628 -613 632 -606
rect 654 -613 658 -606
rect 663 -613 667 -604
rect 672 -613 676 -599
rect 729 -602 734 -601
rect 722 -606 734 -602
rect 693 -614 702 -610
rect 745 -610 748 -593
rect 729 -617 733 -613
rect 744 -614 748 -610
rect 729 -620 736 -617
rect 684 -626 687 -621
rect 684 -633 688 -626
rect 714 -633 718 -626
rect 733 -649 736 -620
rect 637 -662 641 -653
rect 696 -653 706 -649
rect 726 -653 736 -649
rect 646 -665 649 -653
rect 646 -666 655 -665
rect 628 -670 629 -666
rect 637 -669 655 -666
rect 637 -674 641 -669
rect 672 -670 675 -653
rect 703 -660 706 -653
rect 683 -664 685 -660
rect 703 -664 715 -660
rect 703 -665 706 -664
rect 733 -665 736 -653
rect 663 -673 675 -670
rect 663 -674 667 -673
rect 741 -676 744 -614
rect 758 -633 762 -626
rect 774 -635 777 -593
rect 782 -566 789 -563
rect 782 -595 785 -566
rect 831 -572 834 -567
rect 800 -579 804 -572
rect 830 -579 834 -572
rect 782 -599 792 -595
rect 812 -599 822 -595
rect 782 -611 785 -599
rect 812 -606 815 -599
rect 803 -610 815 -606
rect 833 -610 835 -606
rect 812 -611 815 -610
rect 843 -616 846 -599
rect 869 -611 872 -599
rect 877 -608 881 -599
rect 863 -612 872 -611
rect 863 -615 881 -612
rect 843 -619 855 -616
rect 851 -620 855 -619
rect 877 -620 881 -615
rect 889 -616 896 -612
rect 791 -632 795 -631
rect 800 -635 804 -631
rect 821 -632 825 -631
rect 830 -635 834 -631
rect 860 -634 864 -630
rect 886 -634 890 -630
rect 860 -635 890 -634
rect 774 -638 890 -635
rect 899 -641 902 -395
rect 793 -645 816 -641
rect 823 -645 846 -641
rect 853 -645 872 -641
rect 879 -645 902 -641
rect 766 -660 770 -653
rect 753 -664 759 -660
rect 766 -664 776 -660
rect 766 -665 770 -664
rect 758 -676 762 -675
rect 741 -679 762 -676
rect 628 -688 632 -684
rect 654 -688 658 -684
rect 628 -689 658 -688
rect 684 -689 688 -685
rect 693 -686 697 -685
rect 714 -689 718 -685
rect 723 -686 727 -685
rect 741 -689 744 -679
rect 628 -692 744 -689
rect 789 -695 792 -645
rect 813 -649 816 -645
rect 825 -649 828 -645
rect 813 -652 828 -649
rect 843 -649 846 -645
rect 855 -649 858 -645
rect 843 -652 858 -649
rect 869 -649 872 -645
rect 881 -649 884 -645
rect 869 -652 884 -649
rect 453 -741 620 -738
rect 634 -699 639 -695
rect 646 -699 665 -695
rect 672 -699 695 -695
rect 702 -699 725 -695
rect 729 -699 792 -695
rect 634 -703 637 -699
rect 646 -703 649 -699
rect 634 -706 649 -703
rect 660 -703 663 -699
rect 672 -703 675 -699
rect 660 -706 675 -703
rect 690 -703 693 -699
rect 702 -703 705 -699
rect 690 -706 705 -703
rect 453 -751 456 -741
rect 634 -744 637 -706
rect 560 -747 637 -744
rect 383 -755 401 -751
rect 412 -755 419 -751
rect 443 -755 456 -751
rect 483 -755 490 -751
rect 379 -798 383 -773
rect 390 -785 394 -762
rect 397 -760 401 -755
rect 397 -764 402 -760
rect 416 -769 419 -755
rect 397 -779 401 -772
rect 412 -773 415 -769
rect 420 -773 423 -769
rect 397 -782 406 -779
rect 444 -779 448 -762
rect 453 -760 456 -755
rect 453 -764 463 -760
rect 411 -782 448 -779
rect 490 -769 493 -755
rect 452 -785 456 -772
rect 483 -773 493 -769
rect 390 -788 456 -785
rect 429 -790 434 -788
rect 490 -798 493 -773
rect 379 -801 493 -798
rect 310 -807 336 -804
rect 382 -802 387 -801
rect 310 -825 314 -807
rect 395 -809 417 -806
rect 395 -810 399 -809
rect 310 -849 314 -829
rect 303 -852 314 -849
rect 317 -813 395 -810
rect 317 -836 320 -813
rect 416 -810 417 -809
rect 422 -809 479 -806
rect 344 -821 392 -818
rect 323 -831 324 -827
rect 356 -828 360 -821
rect 389 -825 396 -821
rect 403 -825 408 -820
rect 403 -832 407 -825
rect 317 -840 324 -836
rect 303 -861 306 -852
rect 310 -861 314 -859
rect 303 -864 314 -861
rect 310 -879 314 -864
rect 303 -882 314 -879
rect 317 -866 320 -840
rect 345 -848 349 -839
rect 376 -840 383 -836
rect 344 -851 360 -848
rect 323 -861 324 -857
rect 356 -858 360 -851
rect 395 -861 399 -852
rect 317 -870 324 -866
rect 303 -891 306 -882
rect 310 -891 314 -889
rect 303 -894 314 -891
rect 310 -905 314 -894
rect 303 -908 314 -905
rect 317 -896 320 -870
rect 345 -871 349 -869
rect 376 -867 383 -866
rect 376 -870 388 -867
rect 336 -882 356 -879
rect 396 -882 413 -878
rect 336 -887 339 -882
rect 410 -887 413 -882
rect 416 -879 420 -810
rect 454 -879 458 -809
rect 475 -810 479 -809
rect 479 -813 557 -810
rect 466 -825 471 -820
rect 482 -821 530 -818
rect 478 -825 485 -821
rect 467 -832 471 -825
rect 514 -828 518 -821
rect 550 -831 551 -827
rect 491 -840 498 -836
rect 554 -836 557 -813
rect 525 -848 529 -839
rect 550 -840 557 -836
rect 475 -861 479 -852
rect 514 -851 530 -848
rect 514 -858 518 -851
rect 550 -861 551 -857
rect 491 -867 498 -866
rect 486 -870 498 -867
rect 554 -866 557 -840
rect 560 -825 563 -747
rect 560 -849 564 -829
rect 560 -852 571 -849
rect 525 -871 529 -869
rect 550 -870 557 -866
rect 461 -882 478 -878
rect 518 -882 538 -879
rect 335 -891 339 -887
rect 396 -891 405 -887
rect 410 -890 415 -887
rect 461 -887 464 -882
rect 535 -887 538 -882
rect 412 -894 417 -890
rect 424 -894 429 -889
rect 445 -894 450 -889
rect 459 -890 464 -887
rect 457 -894 462 -890
rect 469 -891 478 -887
rect 535 -891 539 -887
rect 317 -900 325 -896
rect 303 -917 306 -908
rect 310 -917 314 -915
rect 303 -920 314 -917
rect 310 -935 314 -920
rect 317 -922 321 -900
rect 340 -905 344 -899
rect 396 -900 403 -896
rect 424 -901 428 -894
rect 340 -908 356 -905
rect 446 -901 450 -894
rect 471 -900 478 -896
rect 554 -896 557 -870
rect 560 -861 564 -859
rect 568 -861 571 -852
rect 560 -864 571 -861
rect 560 -879 564 -864
rect 560 -882 571 -879
rect 530 -905 534 -899
rect 549 -900 557 -896
rect 518 -908 534 -905
rect 340 -913 343 -908
rect 531 -913 534 -908
rect 335 -917 343 -913
rect 347 -917 356 -913
rect 518 -917 527 -913
rect 531 -917 539 -913
rect 317 -926 325 -922
rect 339 -932 343 -925
rect 396 -926 403 -922
rect 406 -929 409 -927
rect 416 -929 420 -921
rect 454 -929 458 -921
rect 471 -926 478 -922
rect 553 -922 557 -900
rect 560 -891 564 -889
rect 568 -891 571 -882
rect 560 -894 571 -891
rect 560 -905 564 -894
rect 560 -908 571 -905
rect 465 -929 468 -927
rect 406 -932 468 -929
rect 531 -932 535 -925
rect 549 -926 557 -922
rect 560 -917 564 -915
rect 568 -917 571 -908
rect 560 -920 571 -917
rect 560 -935 564 -920
rect 310 -938 564 -935
<< m2contact >>
rect 371 -93 377 -87
rect 434 -93 440 -87
rect 371 -119 377 -113
rect 434 -119 440 -113
rect 277 -200 282 -195
rect 351 -152 356 -147
rect 362 -153 368 -148
rect 443 -153 449 -148
rect 455 -152 460 -147
rect 351 -178 356 -173
rect 403 -197 408 -192
rect 455 -178 460 -173
rect 430 -194 435 -189
rect 155 -262 160 -257
rect 224 -251 229 -245
rect 258 -242 264 -236
rect 284 -242 290 -236
rect 199 -262 204 -257
rect 225 -262 230 -257
rect 415 -243 420 -238
rect 684 -222 689 -217
rect 511 -251 516 -246
rect 31 -333 37 -327
rect 57 -333 63 -327
rect 133 -328 138 -323
rect 92 -342 97 -336
rect 91 -353 96 -348
rect 117 -353 122 -348
rect -48 -469 -43 -464
rect -22 -469 -17 -464
rect -108 -490 -102 -484
rect -82 -490 -76 -484
rect -47 -481 -42 -475
rect 25 -397 30 -392
rect 278 -343 283 -338
rect 424 -280 429 -275
rect 300 -366 305 -361
rect 19 -468 24 -463
rect 229 -386 234 -381
rect 300 -385 305 -380
rect -6 -494 -1 -489
rect 8 -517 14 -512
rect -108 -552 -102 -546
rect -82 -552 -76 -546
rect -47 -561 -42 -555
rect -48 -572 -43 -567
rect -22 -572 -17 -567
rect 300 -399 305 -394
rect 479 -326 484 -321
rect 425 -342 430 -337
rect 379 -375 384 -370
rect 257 -410 262 -405
rect 300 -431 305 -426
rect 229 -451 234 -446
rect 245 -450 250 -445
rect 300 -450 305 -445
rect 78 -498 83 -493
rect 39 -508 44 -503
rect 47 -517 53 -512
rect 300 -464 305 -459
rect 257 -475 262 -470
rect 284 -471 289 -466
rect 339 -453 344 -448
rect 363 -481 368 -476
rect 234 -494 239 -489
rect 243 -497 248 -492
rect 259 -523 264 -518
rect 466 -365 471 -360
rect 490 -366 495 -361
rect 634 -296 639 -291
rect 660 -296 665 -291
rect 574 -317 580 -311
rect 600 -317 606 -311
rect 635 -308 640 -302
rect 864 -274 870 -268
rect 748 -286 754 -280
rect 774 -286 780 -280
rect 704 -296 709 -291
rect 809 -295 814 -289
rect 513 -326 518 -321
rect 808 -306 813 -301
rect 834 -306 839 -301
rect 690 -328 695 -323
rect 878 -306 883 -301
rect 490 -393 495 -388
rect 446 -436 451 -431
rect 465 -436 470 -431
rect 479 -436 484 -431
rect 860 -372 865 -367
rect 690 -378 695 -372
rect 742 -379 747 -374
rect 545 -428 550 -423
rect 649 -438 654 -433
rect 439 -457 444 -452
rect 319 -524 324 -519
rect 338 -524 343 -519
rect 352 -524 357 -519
rect 473 -460 479 -454
rect 77 -554 82 -549
rect 252 -547 257 -542
rect 390 -548 395 -543
rect 521 -486 526 -481
rect 603 -466 608 -461
rect 713 -433 718 -428
rect 702 -471 707 -466
rect 539 -496 544 -491
rect 481 -521 487 -516
rect 471 -547 477 -542
rect 489 -536 494 -531
rect 508 -536 513 -531
rect 522 -536 527 -531
rect 531 -538 536 -533
rect 545 -530 550 -525
rect 127 -585 132 -580
rect 422 -561 427 -556
rect 226 -601 231 -596
rect 110 -648 115 -643
rect 183 -612 188 -607
rect 304 -605 309 -600
rect 183 -626 188 -621
rect 238 -626 243 -621
rect 254 -625 259 -620
rect 364 -612 369 -607
rect 184 -645 189 -640
rect 174 -652 180 -646
rect 293 -632 298 -627
rect 309 -631 314 -626
rect 364 -631 369 -626
rect 294 -656 299 -651
rect 208 -662 213 -657
rect 364 -644 369 -639
rect 321 -656 326 -651
rect 384 -592 389 -587
rect 468 -570 473 -565
rect 533 -579 538 -574
rect 403 -648 408 -643
rect 472 -645 477 -640
rect 78 -668 83 -663
rect 208 -690 213 -685
rect 509 -607 514 -602
rect 537 -633 542 -628
rect 731 -508 736 -503
rect 740 -517 745 -512
rect 701 -527 706 -522
rect 571 -605 577 -600
rect 521 -646 527 -641
rect 544 -642 549 -637
rect 583 -658 588 -653
rect 552 -670 557 -665
rect 559 -686 564 -681
rect 235 -757 240 -752
rect 261 -757 266 -752
rect 260 -769 265 -763
rect 294 -778 300 -772
rect 320 -778 326 -772
rect 431 -735 436 -730
rect 462 -735 467 -730
rect 552 -735 557 -730
rect 570 -729 575 -724
rect 584 -729 589 -724
rect 603 -729 608 -724
rect 860 -404 866 -398
rect 800 -469 805 -464
rect 826 -469 831 -464
rect 825 -481 830 -475
rect 784 -494 789 -489
rect 859 -490 865 -484
rect 885 -490 891 -484
rect 769 -503 775 -498
rect 759 -573 764 -568
rect 825 -561 830 -555
rect 859 -552 865 -546
rect 885 -552 891 -546
rect 627 -606 633 -600
rect 653 -606 659 -600
rect 688 -615 693 -609
rect 687 -626 692 -621
rect 713 -626 718 -621
rect 757 -626 762 -621
rect 800 -572 805 -567
rect 826 -572 831 -567
rect 415 -774 420 -769
rect 406 -782 411 -777
rect 382 -807 387 -802
rect 417 -810 422 -805
rect 408 -825 413 -820
rect 383 -841 388 -836
rect 383 -867 388 -862
rect 394 -866 400 -861
rect 486 -841 491 -836
rect 474 -866 480 -861
rect 486 -867 491 -862
rect 403 -901 409 -895
rect 465 -901 471 -895
rect 403 -927 409 -921
rect 465 -927 471 -921
<< metal2 >>
rect 374 -113 377 -93
rect 374 -147 377 -119
rect 434 -113 437 -93
rect 434 -147 437 -119
rect 356 -148 407 -147
rect 356 -150 362 -148
rect 351 -173 354 -152
rect 368 -150 407 -148
rect 434 -148 455 -147
rect 434 -150 443 -148
rect 404 -192 407 -150
rect 449 -150 455 -148
rect 457 -173 460 -152
rect 282 -200 302 -197
rect 227 -239 258 -236
rect 227 -245 230 -239
rect 264 -239 284 -236
rect 229 -251 230 -245
rect 227 -257 230 -251
rect 94 -262 155 -259
rect 160 -262 199 -259
rect 204 -262 225 -259
rect 94 -327 97 -262
rect 37 -330 57 -327
rect 63 -330 97 -327
rect 138 -328 168 -325
rect 91 -336 97 -330
rect 91 -342 92 -336
rect 91 -348 94 -342
rect 96 -353 117 -350
rect 165 -351 168 -328
rect 299 -338 302 -200
rect 430 -223 433 -194
rect 644 -197 714 -192
rect 709 -207 714 -197
rect 709 -212 902 -207
rect 689 -222 902 -217
rect 416 -226 502 -223
rect 416 -238 419 -226
rect 283 -341 302 -338
rect 311 -277 337 -276
rect 311 -279 424 -277
rect 230 -366 300 -363
rect 230 -381 233 -366
rect 21 -392 24 -391
rect 21 -395 25 -392
rect 247 -405 250 -385
rect 300 -394 304 -385
rect 235 -408 257 -405
rect 230 -431 300 -428
rect 230 -446 233 -431
rect -43 -467 -22 -464
rect -17 -467 19 -464
rect -48 -475 -45 -469
rect 247 -470 250 -450
rect 300 -459 304 -450
rect 235 -473 257 -470
rect -48 -481 -47 -475
rect 284 -479 288 -471
rect 227 -481 288 -479
rect -102 -490 -82 -487
rect -48 -487 -45 -481
rect -76 -490 -45 -487
rect 24 -482 288 -481
rect 24 -484 230 -482
rect 24 -491 27 -484
rect 311 -486 314 -279
rect 332 -280 424 -279
rect 425 -337 429 -280
rect 484 -326 485 -321
rect 448 -364 466 -361
rect 384 -373 430 -370
rect 356 -414 408 -411
rect 245 -489 314 -486
rect 321 -452 339 -449
rect -1 -494 27 -491
rect 79 -493 234 -490
rect 24 -504 27 -494
rect 245 -492 248 -489
rect 78 -501 89 -498
rect 24 -507 39 -504
rect 14 -516 47 -513
rect -102 -549 -82 -546
rect -76 -549 -45 -546
rect -48 -555 -45 -549
rect -48 -561 -47 -555
rect -48 -567 -45 -561
rect -43 -572 -22 -569
rect 79 -663 82 -554
rect 86 -589 89 -501
rect 321 -519 324 -452
rect 363 -466 366 -454
rect 404 -456 408 -414
rect 427 -452 430 -373
rect 448 -431 451 -364
rect 490 -378 493 -366
rect 470 -381 493 -378
rect 490 -388 493 -381
rect 499 -388 502 -226
rect 513 -321 516 -251
rect 639 -294 660 -291
rect 665 -294 704 -291
rect 634 -302 637 -296
rect 634 -308 635 -302
rect 580 -317 600 -314
rect 634 -314 637 -308
rect 606 -317 637 -314
rect 512 -326 513 -321
rect 692 -372 695 -328
rect 739 -379 742 -222
rect 808 -232 902 -227
rect 808 -280 811 -232
rect 866 -242 902 -237
rect 866 -268 870 -242
rect 754 -283 774 -280
rect 780 -283 811 -280
rect 808 -289 811 -283
rect 808 -295 809 -289
rect 808 -301 811 -295
rect 813 -306 834 -303
rect 839 -306 878 -303
rect 495 -391 502 -388
rect 862 -398 865 -372
rect 514 -428 545 -425
rect 470 -435 479 -431
rect 427 -455 439 -452
rect 514 -454 517 -428
rect 695 -433 713 -430
rect 479 -457 517 -454
rect 608 -465 675 -462
rect 343 -469 366 -466
rect 363 -476 366 -469
rect 377 -470 524 -467
rect 260 -542 263 -523
rect 343 -523 352 -519
rect 257 -545 263 -542
rect 377 -582 380 -470
rect 521 -481 524 -470
rect 672 -468 675 -465
rect 695 -468 698 -433
rect 672 -471 698 -468
rect 805 -467 826 -464
rect 828 -475 831 -469
rect 830 -481 831 -475
rect 828 -487 831 -481
rect 511 -494 539 -491
rect 511 -516 514 -494
rect 828 -490 859 -487
rect 865 -490 885 -487
rect 736 -506 773 -503
rect 487 -519 514 -516
rect 785 -513 789 -494
rect 745 -516 789 -513
rect 550 -530 705 -527
rect 513 -536 522 -532
rect 395 -547 471 -544
rect 427 -561 471 -558
rect 468 -565 471 -561
rect 132 -585 380 -582
rect 86 -592 384 -589
rect 231 -601 253 -598
rect 304 -599 385 -596
rect 304 -600 309 -599
rect 184 -621 188 -612
rect 238 -621 241 -601
rect 294 -612 364 -609
rect 255 -640 258 -625
rect 294 -627 297 -612
rect 189 -643 258 -640
rect 115 -648 174 -647
rect 110 -650 174 -648
rect 311 -651 314 -631
rect 364 -639 368 -631
rect 382 -643 385 -599
rect 469 -630 472 -570
rect 491 -603 494 -536
rect 757 -534 760 -516
rect 536 -537 760 -534
rect 828 -549 859 -546
rect 828 -555 831 -549
rect 865 -549 885 -546
rect 830 -561 831 -555
rect 828 -567 831 -561
rect 764 -572 800 -569
rect 805 -572 826 -569
rect 533 -586 536 -579
rect 513 -589 536 -586
rect 533 -601 536 -589
rect 491 -606 509 -603
rect 577 -603 627 -600
rect 633 -603 653 -600
rect 659 -603 690 -600
rect 687 -609 690 -603
rect 687 -615 688 -609
rect 687 -621 690 -615
rect 692 -626 713 -623
rect 718 -626 757 -623
rect 469 -633 537 -630
rect 542 -632 556 -629
rect 382 -646 403 -643
rect 477 -641 506 -640
rect 477 -643 521 -641
rect 494 -644 521 -643
rect 299 -654 321 -651
rect 296 -660 299 -656
rect 209 -685 212 -662
rect 296 -663 387 -660
rect 196 -755 235 -752
rect 240 -755 261 -752
rect 263 -763 266 -757
rect 265 -769 266 -763
rect 263 -775 266 -769
rect 263 -778 294 -775
rect 300 -778 320 -775
rect 384 -794 387 -663
rect 436 -735 462 -732
rect 545 -740 548 -642
rect 553 -665 556 -632
rect 588 -657 606 -654
rect 552 -730 555 -670
rect 561 -671 564 -659
rect 561 -674 584 -671
rect 561 -681 564 -674
rect 603 -724 606 -657
rect 575 -728 584 -724
rect 402 -743 548 -740
rect 407 -794 410 -782
rect 384 -797 413 -794
rect 383 -836 386 -807
rect 410 -820 413 -797
rect 417 -805 420 -774
rect 383 -862 386 -841
rect 388 -866 394 -864
rect 400 -866 409 -864
rect 388 -867 409 -866
rect 406 -895 409 -867
rect 465 -866 474 -864
rect 488 -862 491 -841
rect 480 -866 486 -864
rect 465 -867 486 -866
rect 406 -921 409 -901
rect 465 -895 468 -867
rect 465 -921 468 -901
<< m123contact >>
rect 312 -143 317 -138
rect 397 -125 402 -120
rect 409 -125 414 -120
rect 494 -143 499 -138
rect 376 -194 381 -189
rect 252 -216 257 -211
rect 183 -237 188 -232
rect 64 -307 69 -302
rect 164 -301 169 -296
rect 234 -301 239 -296
rect 290 -307 295 -302
rect 388 -232 393 -227
rect 331 -269 336 -264
rect 406 -271 411 -266
rect 245 -385 250 -380
rect 284 -385 289 -380
rect 82 -392 87 -387
rect 230 -410 235 -405
rect -57 -430 -52 -425
rect 284 -450 289 -445
rect 230 -475 235 -470
rect 484 -279 489 -274
rect 323 -288 328 -283
rect 372 -357 377 -352
rect 393 -386 398 -381
rect 351 -414 356 -409
rect -75 -515 -70 -510
rect -75 -526 -70 -521
rect 26 -535 33 -529
rect -6 -547 -1 -542
rect 65 -592 70 -587
rect -57 -611 -52 -606
rect 363 -454 368 -449
rect 338 -469 343 -464
rect 465 -381 470 -376
rect 568 -252 573 -246
rect 625 -257 630 -252
rect 695 -257 700 -252
rect 676 -321 681 -316
rect 607 -342 612 -337
rect 610 -365 615 -360
rect 781 -260 786 -255
rect 850 -281 855 -276
rect 799 -345 804 -340
rect 869 -345 874 -340
rect 465 -420 470 -415
rect 487 -420 492 -415
rect 518 -417 523 -412
rect 603 -417 608 -412
rect 370 -463 375 -458
rect 403 -461 409 -456
rect 835 -430 840 -425
rect 603 -451 608 -446
rect 683 -462 688 -457
rect 338 -508 343 -503
rect 93 -532 98 -527
rect 240 -532 245 -527
rect 267 -549 272 -544
rect 93 -563 98 -558
rect 169 -571 181 -566
rect 435 -484 440 -479
rect 528 -477 533 -472
rect 752 -490 757 -485
rect 518 -503 523 -498
rect 709 -508 714 -503
rect 853 -515 858 -510
rect 384 -563 389 -558
rect 393 -587 398 -582
rect 169 -604 174 -599
rect 253 -601 258 -596
rect 199 -626 204 -621
rect 169 -632 174 -627
rect 348 -631 353 -626
rect 853 -526 858 -521
rect 784 -547 789 -542
rect 508 -552 513 -547
rect 660 -580 665 -575
rect 508 -591 513 -586
rect 531 -606 536 -601
rect 729 -601 734 -596
rect 835 -611 840 -606
rect 254 -656 259 -651
rect 370 -653 375 -648
rect 481 -652 487 -647
rect 327 -713 332 -708
rect 200 -718 205 -713
rect 270 -718 275 -713
rect 191 -757 196 -752
rect 219 -782 224 -777
rect 397 -743 402 -738
rect 560 -659 565 -654
rect 584 -674 589 -669
rect 584 -713 589 -708
rect 678 -665 683 -660
rect 748 -665 753 -660
rect 623 -671 628 -665
rect 490 -755 495 -750
rect 288 -803 293 -798
rect 429 -795 434 -790
rect 461 -825 466 -820
rect 344 -876 349 -871
rect 429 -894 434 -889
rect 440 -894 445 -889
rect 525 -876 530 -871
<< metal3 >>
rect 398 -137 401 -125
rect 312 -138 401 -137
rect 317 -140 401 -138
rect 410 -137 413 -125
rect 410 -138 499 -137
rect 410 -140 494 -138
rect 752 -152 902 -147
rect 743 -163 902 -158
rect 183 -173 902 -168
rect 183 -232 188 -173
rect 695 -183 902 -178
rect 381 -193 392 -189
rect 166 -237 183 -234
rect 237 -215 252 -212
rect 166 -296 169 -237
rect 237 -296 240 -215
rect 389 -227 392 -193
rect 393 -230 498 -227
rect 322 -269 331 -266
rect 322 -283 325 -269
rect 406 -274 411 -271
rect 374 -277 484 -274
rect 322 -286 323 -283
rect 239 -301 240 -296
rect 69 -306 84 -303
rect 81 -387 84 -306
rect 292 -350 295 -307
rect 279 -353 295 -350
rect 279 -357 282 -353
rect 279 -360 287 -357
rect 284 -380 287 -360
rect 81 -392 82 -387
rect 232 -422 235 -410
rect 325 -411 328 -288
rect 374 -352 377 -277
rect 370 -384 393 -381
rect 325 -414 351 -411
rect 495 -415 498 -230
rect 520 -251 568 -247
rect 520 -330 523 -251
rect 695 -252 700 -183
rect 419 -418 465 -415
rect 232 -425 287 -422
rect -58 -430 -57 -425
rect -58 -511 -55 -430
rect 284 -445 287 -425
rect 419 -449 422 -418
rect 492 -418 498 -415
rect 510 -333 523 -330
rect 624 -257 625 -252
rect 850 -193 902 -188
rect 368 -452 422 -449
rect 375 -463 387 -460
rect 409 -461 439 -458
rect 510 -461 513 -333
rect 624 -338 627 -257
rect 695 -316 698 -257
rect 786 -259 801 -256
rect 681 -319 698 -316
rect 612 -341 627 -338
rect 798 -340 801 -259
rect 850 -276 855 -193
rect 855 -281 872 -278
rect 869 -340 872 -281
rect 798 -345 799 -340
rect 606 -365 610 -362
rect 605 -412 608 -365
rect 230 -482 233 -475
rect -70 -514 -55 -511
rect 26 -485 233 -482
rect -70 -525 -55 -522
rect -58 -606 -55 -525
rect 26 -529 29 -485
rect 315 -506 338 -503
rect -6 -535 26 -531
rect 245 -532 270 -529
rect -6 -542 -2 -535
rect 93 -558 96 -532
rect 267 -544 270 -532
rect 315 -567 318 -506
rect 384 -558 387 -463
rect 436 -479 439 -461
rect 477 -464 513 -461
rect 477 -528 480 -464
rect 518 -474 521 -417
rect 603 -446 606 -417
rect 840 -430 841 -425
rect 518 -477 528 -474
rect 683 -474 686 -462
rect 607 -477 713 -474
rect 518 -487 521 -477
rect 607 -487 610 -477
rect 518 -490 610 -487
rect 518 -498 521 -490
rect 710 -503 713 -477
rect 757 -490 758 -485
rect 755 -528 758 -490
rect 838 -511 841 -430
rect 838 -514 853 -511
rect 838 -525 853 -522
rect 397 -531 480 -528
rect 552 -531 789 -528
rect 397 -567 400 -531
rect 315 -570 400 -567
rect 485 -552 508 -549
rect 173 -586 176 -571
rect 170 -587 176 -586
rect 70 -589 176 -587
rect 70 -590 173 -589
rect 170 -599 173 -590
rect 300 -596 351 -593
rect 300 -598 303 -596
rect 258 -601 303 -598
rect -58 -611 -57 -606
rect 170 -653 173 -632
rect 201 -646 204 -626
rect 348 -626 351 -596
rect 201 -649 208 -646
rect 170 -656 254 -653
rect 170 -752 173 -656
rect 372 -658 375 -653
rect 372 -661 389 -658
rect 327 -708 332 -704
rect 275 -718 276 -713
rect 170 -755 191 -752
rect 202 -777 205 -718
rect 202 -780 219 -777
rect 219 -805 224 -782
rect 273 -799 276 -718
rect 386 -794 389 -661
rect 394 -741 397 -587
rect 485 -640 488 -552
rect 552 -601 555 -531
rect 785 -542 789 -531
rect 665 -579 680 -576
rect 536 -604 555 -601
rect 485 -643 501 -640
rect 498 -647 501 -643
rect 487 -652 494 -649
rect 498 -650 563 -647
rect 491 -750 494 -652
rect 560 -654 563 -650
rect 677 -660 680 -579
rect 734 -601 748 -598
rect 748 -660 751 -603
rect 838 -606 841 -525
rect 840 -611 841 -606
rect 677 -665 678 -660
rect 609 -670 623 -666
rect 609 -708 612 -670
rect 589 -711 612 -708
rect 386 -795 429 -794
rect 434 -795 464 -794
rect 386 -797 464 -795
rect 273 -802 288 -799
rect 461 -820 464 -797
rect 349 -876 433 -874
rect 344 -877 433 -876
rect 430 -889 433 -877
rect 441 -876 525 -874
rect 441 -877 530 -876
rect 441 -889 444 -877
<< m234contact >>
rect 639 -197 644 -192
rect 19 -391 24 -386
rect 164 -356 169 -351
rect 485 -326 490 -321
rect 507 -326 512 -321
rect 601 -365 606 -360
<< m4contact >>
rect 747 -152 752 -147
rect 738 -163 743 -158
rect 365 -385 370 -380
rect 208 -649 213 -644
rect 327 -704 332 -699
rect 748 -603 753 -598
rect 219 -810 224 -805
<< metal4 >>
rect 159 -196 639 -192
rect 159 -252 163 -196
rect 740 -208 743 -163
rect 133 -256 163 -252
rect 375 -211 743 -208
rect 133 -296 137 -256
rect 20 -300 137 -296
rect 20 -386 24 -300
rect 169 -355 317 -352
rect 314 -380 317 -355
rect 314 -383 365 -380
rect 213 -649 249 -646
rect 246 -668 249 -649
rect 246 -671 332 -668
rect 327 -699 332 -671
rect 375 -807 378 -211
rect 490 -326 507 -323
rect 507 -362 510 -326
rect 507 -365 601 -362
rect 749 -598 752 -152
rect 224 -810 378 -807
<< labels >>
rlabel metal3 486 -563 486 -563 1 node31
rlabel metal3 342 -595 346 -594 1 node21
rlabel metal3 273 -424 277 -423 1 node11
rlabel metal3 434 -417 435 -416 1 node01
rlabel metal1 474 -489 476 -484 1 Pout_bar
rlabel metal1 541 -499 541 -499 1 node34
rlabel metal1 567 -436 567 -436 1 node35
rlabel metal1 651 -441 651 -441 1 node33
rlabel metal1 671 -480 671 -480 1 node32
rlabel metal1 559 -708 559 -708 1 C3
rlabel metal1 332 -327 332 -327 1 C1
rlabel metal1 490 -605 490 -605 1 node25
rlabel metal1 487 -689 487 -689 1 node23
rlabel metal1 429 -579 429 -579 1 node24
rlabel metal1 447 -709 447 -709 1 node22
rlabel metal1 113 -641 113 -641 1 C2
rlabel metal1 133 -579 133 -579 1 node13
rlabel metal1 216 -586 216 -586 1 node15
rlabel metal1 243 -526 243 -526 1 node14
rlabel metal1 112 -545 112 -545 1 node12
rlabel metal1 367 -339 367 -339 1 node02
rlabel metal1 546 -373 548 -371 1 node36
rlabel metal1 670 -396 672 -393 1 Gout_bar
rlabel metal1 710 -470 712 -468 1 G3_bar
rlabel metal1 710 -525 712 -523 1 P3_bar
rlabel metal1 398 -749 400 -747 1 P2_bar
rlabel metal1 453 -749 455 -747 1 G2_bar
rlabel metal1 72 -552 74 -550 1 G1_bar
rlabel metal1 72 -497 74 -495 1 P1_bar
rlabel metal1 426 -273 428 -271 1 P0_bar
rlabel metal1 371 -273 373 -271 1 G0_bar
rlabel metal1 419 -511 421 -509 1 C0_bar
rlabel metal1 890 -615 891 -613 1 A3
rlabel metal1 -108 -615 -107 -613 1 A1
rlabel metal1 -108 -423 -107 -421 1 B1
rlabel metal1 308 -88 310 -87 5 A0
rlabel metal3 866 -183 902 -178 1 S0
rlabel metal3 866 -163 902 -158 1 S2
rlabel metal3 866 -152 902 -147 1 S3
rlabel metal3 866 -193 902 -188 1 Cout
rlabel metal2 866 -222 902 -217 1 clk
rlabel metal2 866 -232 902 -227 1 vdd
rlabel metal2 866 -242 902 -237 1 gnd
rlabel metal1 891 -423 894 -421 1 B3
rlabel metal2 866 -212 902 -207 1 C0
rlabel metal1 501 -88 503 -87 5 B0
rlabel metal1 340 -930 342 -927 1 B2
rlabel metal1 532 -930 534 -927 1 A2
rlabel metal3 866 -173 902 -168 1 S1
rlabel metal3 389 -216 392 -212 1 A0_after
rlabel metal2 430 -216 433 -212 1 B0_after
rlabel metal3 13 -535 19 -531 1 A1_after
rlabel metal2 14 -494 19 -491 1 B1_after
rlabel metal3 461 -805 464 -801 1 A2_after
rlabel metal2 410 -805 413 -801 1 B2_after
rlabel metal3 764 -531 769 -528 1 A3_after
rlabel metal2 764 -516 769 -513 1 B3_after
rlabel metal3 553 -251 561 -247 1 S0_before
rlabel metal3 292 -320 295 -315 1 S1_before
rlabel metal4 328 -694 331 -689 1 S2_before
rlabel metal3 609 -676 612 -671 1 S3_before
rlabel metal1 726 -350 733 -346 1 Cout_before
rlabel metal2 165 -337 168 -330 1 C0_after
<< end >>
