magic
tech scmos
timestamp 1731177396
<< nwell >>
rect -1 -38 49 -6
<< ntransistor >>
rect 10 -72 12 -52
rect 20 -72 22 -52
rect 36 -54 38 -44
<< ptransistor >>
rect 10 -32 12 -12
rect 20 -32 22 -12
rect 36 -32 38 -12
<< ndiffusion >>
rect 31 -50 36 -44
rect 5 -68 10 -52
rect 9 -72 10 -68
rect 12 -72 20 -52
rect 22 -56 23 -52
rect 35 -54 36 -50
rect 38 -48 39 -44
rect 38 -54 43 -48
rect 22 -72 27 -56
<< pdiffusion >>
rect 9 -16 10 -12
rect 5 -32 10 -16
rect 12 -28 20 -12
rect 12 -32 14 -28
rect 18 -32 20 -28
rect 22 -16 23 -12
rect 22 -32 27 -16
rect 35 -16 36 -12
rect 31 -32 36 -16
rect 38 -28 43 -12
rect 38 -32 39 -28
<< ndcontact >>
rect 5 -72 9 -68
rect 23 -56 27 -52
rect 31 -54 35 -50
rect 39 -48 43 -44
<< pdcontact >>
rect 5 -16 9 -12
rect 14 -32 18 -28
rect 23 -16 27 -12
rect 31 -16 35 -12
rect 39 -32 43 -28
<< polysilicon >>
rect 10 -12 12 -8
rect 20 -12 22 -8
rect 36 -12 38 -8
rect 10 -52 12 -32
rect 20 -52 22 -32
rect 36 -44 38 -32
rect 36 -58 38 -54
rect 10 -75 12 -72
rect 20 -75 22 -72
<< polycontact >>
rect 6 -43 10 -39
rect 16 -51 20 -47
rect 32 -43 36 -39
<< metal1 >>
rect 5 -5 35 -2
rect 5 -12 9 -5
rect 23 -12 27 -5
rect 31 -12 35 -5
rect 14 -39 18 -32
rect 39 -39 43 -32
rect -1 -43 6 -39
rect 14 -43 32 -39
rect 39 -43 49 -39
rect -1 -51 16 -47
rect 23 -52 27 -43
rect 39 -44 43 -43
rect 5 -76 9 -72
rect 31 -76 35 -54
rect 5 -79 35 -76
<< labels >>
rlabel metal1 15 -4 17 -3 5 vdd
rlabel metal1 1 -41 3 -40 3 a
rlabel metal1 3 -50 4 -48 3 b
rlabel metal1 6 -74 8 -73 1 gnd
rlabel metal1 46 -42 48 -40 7 out
<< end >>
