* SPICE3 file created from and_layout.ext - technology: scmos

.include TSMC_180nm.txt
.param vdd=1.8
.param LAMBDA=0.09u
.global vdd gnd
.option scale=0.09u

M1000 a_12_n32# a vdd w_n1_n38# CMOSP w=20 l=2
+  ad=160 pd=56 as=300 ps=150
M1001 a_12_n72# a gnd Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=150 ps=80
M1002 vdd b a_12_n32# w_n1_n38# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_12_n32# b a_12_n72# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1004 out a_12_n32# vdd w_n1_n38# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1005 out a_12_n32# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 a_12_n32# gnd 0.09fF
C1 b a 0.21fF
C2 a_12_n32# w_n1_n38# 0.09fF
C3 out w_n1_n38# 0.02fF
C4 a_12_n32# out 0.05fF
C5 b w_n1_n38# 0.07fF
C6 b a_12_n32# 0.19fF
C7 w_n1_n38# a 0.07fF
C8 a_12_n32# a 0.04fF
C9 vdd w_n1_n38# 0.07fF
C10 gnd Gnd 0.01fF
C11 out Gnd 0.04fF
C12 vdd Gnd 0.08fF
C13 a_12_n32# Gnd 0.19fF
C14 b Gnd 0.19fF
C15 a Gnd 0.16fF
C16 w_n1_n38# Gnd 1.61fF

Vdd vdd gnd dc 1.8
* trise = tfall = 5% of T_on
Va  a  gnd pulse 1.8 0 5n 100ps  100ps  10ns 20ns
Vb  b  gnd pulse 1.8 0 0  100ps  100ps  20ns 40ns
* .ic v(out) = 0
.tran 1ps 200ns 1ps
* CL out gnd 50f

* clk - out propagation delay
.measure tran t_rise TRIG V(a) VAL='0.9' FALL=1 TARG V(out) VAL='0.9' RISE=1
.measure tran t_fall TRIG V(a) VAL='0.9' RISE=2 TARG V(out) VAL='0.9' FALL=1
.measure tran prop_delay param ='(t_rise + t_fall)/2'

* 20lambda: 304p, 245p, 275p
* saturates around 90p

.control
set hcopypscolor = 1
set color0 = white
set color1 = black

run
set curplottitle= "M P Samartha-2023102038"
plot a+4, b+2, out
.endc





