magic
tech scmos
timestamp 1731158097
<< nwell >>
rect 0 0 34 32
<< ntransistor >>
rect 11 -34 13 -14
rect 21 -34 23 -14
<< ptransistor >>
rect 11 6 13 26
rect 21 6 23 26
<< ndiffusion >>
rect 6 -30 11 -14
rect 10 -34 11 -30
rect 13 -34 21 -14
rect 23 -18 24 -14
rect 23 -34 28 -18
<< pdiffusion >>
rect 10 22 11 26
rect 6 6 11 22
rect 13 10 21 26
rect 13 6 15 10
rect 19 6 21 10
rect 23 22 24 26
rect 23 6 28 22
<< ndcontact >>
rect 6 -34 10 -30
rect 24 -18 28 -14
<< pdcontact >>
rect 6 22 10 26
rect 15 6 19 10
rect 24 22 28 26
<< polysilicon >>
rect 11 26 13 30
rect 21 26 23 30
rect 11 -14 13 6
rect 21 -14 23 6
rect 11 -37 13 -34
rect 21 -37 23 -34
<< polycontact >>
rect 7 -5 11 -1
rect 17 -13 21 -9
<< metal1 >>
rect 6 33 28 36
rect 6 26 10 33
rect 24 26 28 33
rect 15 -1 19 6
rect 0 -5 7 -1
rect 15 -5 34 -1
rect 0 -13 17 -9
rect 24 -14 28 -5
rect 6 -37 10 -34
<< labels >>
rlabel metal1 16 34 18 35 5 vdd
rlabel metal1 2 -3 4 -2 3 a
rlabel metal1 4 -12 5 -10 3 b
rlabel metal1 30 -4 32 -2 1 out
rlabel metal1 7 -36 9 -35 1 gnd
<< end >>
