magic
tech scmos
timestamp 1731237221
<< error_s >>
rect 27 20 30 52
<< nwell >>
rect -42 -17 -18 15
<< ntransistor >>
rect -31 -33 -29 -23
<< ptransistor >>
rect -31 -11 -29 9
<< ndiffusion >>
rect -36 -29 -31 -23
rect -32 -33 -31 -29
rect -29 -27 -28 -23
rect -29 -33 -24 -27
<< pdiffusion >>
rect -32 5 -31 9
rect -36 -11 -31 5
rect -29 -7 -24 9
rect -29 -11 -28 -7
<< ndcontact >>
rect -36 -33 -32 -29
rect -28 -27 -24 -23
<< pdcontact >>
rect -36 5 -32 9
rect -28 -11 -24 -7
<< polysilicon >>
rect -31 9 -29 13
rect -31 -23 -29 -11
rect -31 -37 -29 -33
<< polycontact >>
rect -35 -22 -31 -18
<< metal1 >>
rect -36 9 -32 19
rect -28 -18 -24 -11
rect -42 -22 -35 -18
rect -28 -22 -18 -18
rect -28 -23 -24 -22
rect -36 -37 -32 -33
use not_layout  not_layout_1
timestamp 1731149861
transform 1 0 27 0 1 20
box 0 -20 24 36
use not_layout  not_layout_0
timestamp 1731149861
transform 1 0 0 0 1 20
box 0 -20 24 36
<< labels >>
rlabel metal1 -41 -21 -39 -19 3 in
rlabel metal1 -35 -36 -33 -34 1 gnd
rlabel metal1 -21 -21 -19 -19 7 out
rlabel metal1 -35 16 -33 18 5 vdd
<< end >>
