magic
tech scmos
timestamp 1731356613
<< nwell >>
rect -58 235 -26 269
rect 42 235 94 269
rect -64 192 -30 224
rect -23 173 29 225
rect -230 91 -198 134
rect 67 128 99 171
rect 122 147 154 171
rect -175 91 -143 115
rect -479 20 -455 52
rect -353 24 -319 76
rect -230 37 -198 80
rect -59 61 -35 93
rect 155 88 207 140
rect 221 128 253 162
rect 221 84 273 119
rect -175 37 -143 61
rect -479 -35 -436 -3
rect -279 -36 -227 16
rect -214 -18 -162 16
rect -78 6 -35 38
rect 3 3 27 35
rect 175 27 207 77
rect 221 43 253 77
rect 313 44 347 76
rect 156 -16 208 18
rect 221 -16 273 36
rect -353 -76 -319 -44
rect -259 -77 -227 -43
rect -213 -77 -181 -27
rect 313 -76 347 -24
rect -279 -136 -227 -84
rect 3 -130 37 -78
rect 46 -129 96 -97
rect 3 -195 55 -143
rect 62 -175 96 -143
rect 103 -195 155 -143
rect -58 -269 -6 -235
rect 62 -269 94 -235
<< ntransistor >>
rect -12 256 8 258
rect 19 256 29 258
rect -12 246 8 248
rect 19 246 29 248
rect -53 158 -51 178
rect -43 158 -41 178
rect -12 157 -10 167
rect 6 150 8 160
rect 16 150 18 160
rect 51 158 61 160
rect 105 158 115 160
rect 267 149 287 151
rect 51 139 61 141
rect 267 139 287 141
rect 139 127 149 129
rect -246 121 -236 123
rect 132 109 142 111
rect -246 102 -236 104
rect -192 102 -182 104
rect 286 105 296 107
rect 132 99 142 101
rect 286 95 296 97
rect -246 67 -236 69
rect 159 64 169 66
rect 267 64 287 66
rect -246 48 -236 50
rect -192 48 -182 50
rect -48 44 -46 54
rect 267 54 287 56
rect 141 48 161 50
rect 141 38 161 40
rect -468 3 -466 13
rect -342 1 -340 11
rect -332 1 -330 11
rect -302 3 -292 5
rect -149 3 -139 5
rect 279 23 289 25
rect -302 -7 -292 -5
rect -149 -7 -139 -5
rect -342 -30 -340 -10
rect -332 -30 -330 -10
rect -67 -10 -65 0
rect -48 -10 -46 0
rect 324 10 326 30
rect 334 10 336 30
rect 133 5 143 7
rect 286 5 296 7
rect 14 -13 16 -3
rect 133 -5 143 -3
rect 286 -5 296 -3
rect 324 -11 326 -1
rect 334 -11 336 -1
rect -295 -25 -285 -23
rect -468 -51 -466 -41
rect -449 -51 -447 -41
rect -167 -40 -147 -38
rect -167 -50 -147 -48
rect -293 -56 -273 -54
rect -293 -66 -273 -64
rect -175 -66 -165 -64
rect 14 -65 16 -55
rect 24 -65 26 -55
rect 57 -83 59 -63
rect 67 -83 69 -63
rect -302 -97 -292 -95
rect -302 -107 -292 -105
rect -295 -125 -285 -123
rect 83 -91 85 -81
rect 14 -218 16 -208
rect 24 -218 26 -208
rect 42 -211 44 -201
rect 73 -209 75 -189
rect 83 -209 85 -189
rect 114 -218 116 -208
rect 124 -218 126 -208
rect 142 -211 144 -201
rect 7 -248 17 -246
rect 28 -248 48 -246
rect 7 -258 17 -256
rect 28 -258 48 -256
<< ptransistor >>
rect -52 256 -32 258
rect 48 256 88 258
rect -52 246 -32 248
rect 48 246 88 248
rect -53 198 -51 218
rect -43 198 -41 218
rect -12 179 -10 199
rect 6 179 8 219
rect 16 179 18 219
rect 73 158 93 160
rect 128 158 148 160
rect 227 149 247 151
rect 73 139 93 141
rect 227 139 247 141
rect 161 127 181 129
rect -224 121 -204 123
rect 161 109 201 111
rect -224 102 -204 104
rect -169 102 -149 104
rect 227 105 267 107
rect 161 99 201 101
rect 227 95 267 97
rect -468 26 -466 46
rect -342 30 -340 70
rect -332 30 -330 70
rect -224 67 -204 69
rect -48 67 -46 87
rect 181 64 201 66
rect 227 64 247 66
rect -224 48 -204 50
rect -169 48 -149 50
rect 227 54 247 56
rect 181 48 201 50
rect 324 50 326 70
rect 334 50 336 70
rect 181 38 201 40
rect -67 12 -65 32
rect -48 12 -46 32
rect -273 3 -233 5
rect -208 3 -168 5
rect 14 9 16 29
rect 247 23 267 25
rect -273 -7 -233 -5
rect -208 -7 -168 -5
rect -468 -29 -466 -9
rect -449 -29 -447 -9
rect 162 5 202 7
rect 227 5 267 7
rect 162 -5 202 -3
rect 227 -5 267 -3
rect -273 -25 -253 -23
rect -207 -40 -187 -38
rect -342 -70 -340 -50
rect -332 -70 -330 -50
rect -207 -50 -187 -48
rect -253 -56 -233 -54
rect -253 -66 -233 -64
rect -207 -66 -187 -64
rect 324 -70 326 -30
rect 334 -70 336 -30
rect -273 -97 -233 -95
rect -273 -107 -233 -105
rect -273 -125 -253 -123
rect 14 -124 16 -84
rect 24 -124 26 -84
rect 57 -123 59 -103
rect 67 -123 69 -103
rect 83 -123 85 -103
rect 14 -189 16 -149
rect 24 -189 26 -149
rect 73 -169 75 -149
rect 83 -169 85 -149
rect 42 -189 44 -169
rect 114 -189 116 -149
rect 124 -189 126 -149
rect 142 -189 144 -169
rect -52 -248 -12 -246
rect 68 -248 88 -246
rect -52 -258 -12 -256
rect 68 -258 88 -256
<< ndiffusion >>
rect -12 259 4 263
rect -12 258 8 259
rect 23 259 29 263
rect 19 258 29 259
rect -12 248 8 256
rect 19 254 29 256
rect 19 250 25 254
rect 19 248 29 250
rect -12 245 8 246
rect -8 241 8 245
rect 19 245 29 246
rect 23 241 29 245
rect -54 174 -53 178
rect -58 158 -53 174
rect -51 158 -43 178
rect -41 162 -36 178
rect -41 158 -40 162
rect -13 163 -12 167
rect -17 157 -12 163
rect -10 161 -5 167
rect -10 157 -9 161
rect 55 161 61 165
rect 51 160 61 161
rect 109 161 115 165
rect 105 160 115 161
rect 1 154 6 160
rect 5 150 6 154
rect 8 156 10 160
rect 14 156 16 160
rect 8 150 16 156
rect 18 154 23 160
rect 18 150 19 154
rect 51 157 61 158
rect 51 153 57 157
rect 105 157 115 158
rect 105 153 111 157
rect 271 152 287 156
rect 267 151 287 152
rect 51 142 57 146
rect 51 141 61 142
rect 267 141 287 149
rect 51 138 61 139
rect 51 134 57 138
rect 267 138 287 139
rect 267 134 283 138
rect 139 130 145 134
rect 139 129 149 130
rect -246 124 -240 128
rect -246 123 -236 124
rect 139 126 149 127
rect 143 122 149 126
rect -246 120 -236 121
rect -246 116 -240 120
rect 136 112 142 116
rect 132 111 142 112
rect -246 105 -240 109
rect -246 104 -236 105
rect -192 105 -186 109
rect -192 104 -182 105
rect 132 107 142 109
rect 132 103 138 107
rect -246 101 -236 102
rect -242 97 -236 101
rect -192 101 -182 102
rect -188 97 -182 101
rect 132 101 142 103
rect 286 108 292 112
rect 286 107 296 108
rect 132 98 142 99
rect 136 94 142 98
rect 286 103 296 105
rect 290 99 296 103
rect 286 97 296 99
rect 286 94 296 95
rect 286 90 292 94
rect -246 70 -240 74
rect -246 69 -236 70
rect 159 67 165 71
rect -246 66 -236 67
rect -246 62 -240 66
rect -246 51 -240 55
rect -246 50 -236 51
rect -192 51 -186 55
rect -192 50 -182 51
rect 159 66 169 67
rect 271 67 287 71
rect 267 66 287 67
rect 159 63 169 64
rect 163 59 169 63
rect 267 56 287 64
rect -49 50 -48 54
rect -246 47 -236 48
rect -242 43 -236 47
rect -192 47 -182 48
rect -188 43 -182 47
rect -53 44 -48 50
rect -46 48 -41 54
rect 141 51 157 55
rect 141 50 161 51
rect 267 53 287 54
rect 267 49 283 53
rect -46 44 -45 48
rect 141 40 161 48
rect 141 37 161 38
rect 145 33 161 37
rect -473 7 -468 13
rect -469 3 -468 7
rect -466 9 -465 13
rect -466 3 -461 9
rect -347 5 -342 11
rect -343 1 -342 5
rect -340 7 -338 11
rect -334 7 -332 11
rect -340 1 -332 7
rect -330 5 -325 11
rect -298 6 -292 10
rect -302 5 -292 6
rect -149 6 -143 10
rect -149 5 -139 6
rect -330 1 -329 5
rect -302 1 -292 3
rect -302 -3 -296 1
rect -302 -5 -292 -3
rect -149 1 -139 3
rect -145 -3 -139 1
rect 283 26 289 30
rect 279 25 289 26
rect 323 26 324 30
rect 279 22 289 23
rect 279 18 285 22
rect -149 -5 -139 -3
rect -68 -4 -67 0
rect -302 -8 -292 -7
rect -343 -14 -342 -10
rect -347 -30 -342 -14
rect -340 -30 -332 -10
rect -330 -26 -325 -10
rect -298 -12 -292 -8
rect -149 -8 -139 -7
rect -149 -12 -143 -8
rect -72 -10 -67 -4
rect -65 -4 -64 0
rect -65 -10 -60 -4
rect -49 -4 -48 0
rect -53 -10 -48 -4
rect -46 -6 -41 0
rect 137 8 143 12
rect 133 7 143 8
rect 286 8 292 12
rect 319 10 324 26
rect 326 10 334 30
rect 336 14 341 30
rect 336 10 337 14
rect 286 7 296 8
rect 133 3 143 5
rect 133 -1 139 3
rect 133 -3 143 -1
rect 286 3 296 5
rect 290 -1 296 3
rect 286 -3 296 -1
rect -46 -10 -45 -6
rect 9 -9 14 -3
rect 13 -13 14 -9
rect 16 -7 17 -3
rect 323 -5 324 -1
rect 16 -13 21 -7
rect 133 -6 143 -5
rect 137 -10 143 -6
rect 286 -6 296 -5
rect 286 -10 292 -6
rect 319 -11 324 -5
rect 326 -7 334 -1
rect 326 -11 328 -7
rect 332 -11 334 -7
rect 336 -5 337 -1
rect 336 -11 341 -5
rect -291 -22 -285 -18
rect -295 -23 -285 -22
rect -330 -30 -329 -26
rect -295 -26 -285 -25
rect -295 -30 -289 -26
rect -473 -47 -468 -41
rect -469 -51 -468 -47
rect -466 -45 -465 -41
rect -466 -51 -461 -45
rect -450 -45 -449 -41
rect -454 -51 -449 -45
rect -447 -45 -446 -41
rect -447 -51 -442 -45
rect -167 -37 -151 -33
rect -167 -38 -147 -37
rect -167 -48 -147 -40
rect -289 -53 -273 -49
rect -293 -54 -273 -53
rect -167 -51 -147 -50
rect -163 -55 -147 -51
rect -293 -64 -273 -56
rect 13 -59 14 -55
rect -175 -63 -169 -59
rect -175 -64 -165 -63
rect 9 -65 14 -59
rect 16 -61 24 -55
rect 16 -65 18 -61
rect 22 -65 24 -61
rect 26 -59 27 -55
rect 26 -65 31 -59
rect -293 -67 -273 -66
rect -293 -71 -277 -67
rect -175 -67 -165 -66
rect -171 -71 -165 -67
rect 56 -67 57 -63
rect 52 -83 57 -67
rect 59 -83 67 -63
rect 69 -79 74 -63
rect 69 -83 70 -79
rect -298 -94 -292 -90
rect -302 -95 -292 -94
rect -302 -99 -292 -97
rect -302 -103 -296 -99
rect -302 -105 -292 -103
rect -302 -108 -292 -107
rect -298 -112 -292 -108
rect -291 -122 -285 -118
rect -295 -123 -285 -122
rect 82 -85 83 -81
rect 78 -91 83 -85
rect 85 -87 90 -81
rect 85 -91 86 -87
rect -295 -126 -285 -125
rect -295 -130 -289 -126
rect 37 -207 42 -201
rect 9 -214 14 -208
rect 13 -218 14 -214
rect 16 -212 18 -208
rect 22 -212 24 -208
rect 16 -218 24 -212
rect 26 -214 31 -208
rect 41 -211 42 -207
rect 44 -205 45 -201
rect 44 -211 49 -205
rect 68 -205 73 -189
rect 72 -209 73 -205
rect 75 -209 83 -189
rect 85 -193 86 -189
rect 85 -209 90 -193
rect 137 -207 142 -201
rect 26 -218 27 -214
rect 109 -214 114 -208
rect 113 -218 114 -214
rect 116 -212 118 -208
rect 122 -212 124 -208
rect 116 -218 124 -212
rect 126 -214 131 -208
rect 141 -211 142 -207
rect 144 -205 145 -201
rect 144 -211 149 -205
rect 126 -218 127 -214
rect 7 -245 13 -241
rect 7 -246 17 -245
rect 28 -245 44 -241
rect 28 -246 48 -245
rect 7 -250 17 -248
rect 11 -254 17 -250
rect 7 -256 17 -254
rect 28 -256 48 -248
rect 7 -259 17 -258
rect 7 -263 13 -259
rect 28 -259 48 -258
rect 32 -263 48 -259
<< pdiffusion >>
rect -48 259 -32 263
rect -52 258 -32 259
rect 48 259 84 263
rect 48 258 88 259
rect -52 254 -32 256
rect -52 250 -36 254
rect -52 248 -32 250
rect 48 248 88 256
rect -52 245 -32 246
rect -48 241 -32 245
rect 48 245 88 246
rect 52 241 88 245
rect -54 214 -53 218
rect -58 198 -53 214
rect -51 202 -43 218
rect -51 198 -49 202
rect -45 198 -43 202
rect -41 214 -40 218
rect -41 198 -36 214
rect -17 183 -12 199
rect -13 179 -12 183
rect -10 195 -9 199
rect -10 179 -5 195
rect 1 183 6 219
rect 5 179 6 183
rect 8 179 16 219
rect 18 215 19 219
rect 18 179 23 215
rect 73 161 89 165
rect 73 160 93 161
rect 128 161 144 165
rect 128 160 148 161
rect 73 157 93 158
rect 77 153 93 157
rect 128 157 148 158
rect 132 153 148 157
rect 231 152 247 156
rect 227 151 247 152
rect 227 147 247 149
rect 77 142 93 146
rect 73 141 93 142
rect 227 143 243 147
rect 227 141 247 143
rect 73 138 93 139
rect 77 134 93 138
rect 227 138 247 139
rect 231 134 247 138
rect 165 130 181 134
rect 161 129 181 130
rect -220 124 -204 128
rect -224 123 -204 124
rect 161 126 181 127
rect 161 122 177 126
rect -224 120 -204 121
rect -220 116 -204 120
rect 165 112 201 116
rect 161 111 201 112
rect -220 105 -204 109
rect -224 104 -204 105
rect -165 105 -149 109
rect -169 104 -149 105
rect -224 101 -204 102
rect -224 97 -208 101
rect -169 101 -149 102
rect 161 101 201 109
rect 227 108 263 112
rect 227 107 267 108
rect -169 97 -153 101
rect 161 98 201 99
rect 161 94 197 98
rect 227 97 267 105
rect 227 94 267 95
rect 231 90 267 94
rect -343 66 -342 70
rect -469 42 -468 46
rect -473 26 -468 42
rect -466 30 -461 46
rect -347 30 -342 66
rect -340 30 -332 70
rect -330 34 -325 70
rect -220 70 -204 74
rect -224 69 -204 70
rect -53 71 -48 87
rect -49 67 -48 71
rect -46 83 -45 87
rect -46 67 -41 83
rect -224 66 -204 67
rect -220 62 -204 66
rect -220 51 -204 55
rect -224 50 -204 51
rect -165 51 -149 55
rect 185 67 201 71
rect 181 66 201 67
rect 231 67 247 71
rect 227 66 247 67
rect 323 66 324 70
rect 181 63 201 64
rect 181 59 197 63
rect 227 62 247 64
rect 227 58 243 62
rect 227 56 247 58
rect -169 50 -149 51
rect -224 47 -204 48
rect -224 43 -208 47
rect -169 47 -149 48
rect -169 43 -153 47
rect 181 51 197 55
rect 181 50 201 51
rect 227 53 247 54
rect 231 49 247 53
rect 319 50 324 66
rect 326 54 334 70
rect 326 50 328 54
rect 332 50 334 54
rect 336 66 337 70
rect 336 50 341 66
rect -330 30 -329 34
rect 181 46 201 48
rect 185 42 201 46
rect 181 40 201 42
rect 181 37 201 38
rect 181 33 197 37
rect -466 26 -465 30
rect -72 16 -67 32
rect -68 12 -67 16
rect -65 16 -60 32
rect -65 12 -64 16
rect -53 16 -48 32
rect -49 12 -48 16
rect -46 28 -45 32
rect -46 12 -41 28
rect 13 25 14 29
rect -273 6 -237 10
rect -273 5 -233 6
rect -204 6 -168 10
rect -208 5 -168 6
rect -273 -5 -233 3
rect -208 -5 -168 3
rect 9 9 14 25
rect 16 13 21 29
rect 247 26 263 30
rect 247 25 267 26
rect 247 22 267 23
rect 251 18 267 22
rect 16 9 17 13
rect -469 -13 -468 -9
rect -473 -29 -468 -13
rect -466 -25 -461 -9
rect -466 -29 -465 -25
rect -454 -25 -449 -9
rect -450 -29 -449 -25
rect -447 -25 -442 -9
rect -447 -29 -446 -25
rect -273 -8 -233 -7
rect -269 -12 -233 -8
rect -208 -8 -168 -7
rect -208 -12 -172 -8
rect 166 8 202 12
rect 162 7 202 8
rect 227 8 263 12
rect 227 7 267 8
rect 162 -3 202 5
rect 227 -3 267 5
rect 162 -6 202 -5
rect 162 -10 198 -6
rect 227 -6 267 -5
rect 231 -10 267 -6
rect -273 -22 -257 -18
rect -273 -23 -253 -22
rect -273 -26 -253 -25
rect -269 -30 -253 -26
rect -203 -37 -187 -33
rect -207 -38 -187 -37
rect 323 -34 324 -30
rect -207 -42 -187 -40
rect -207 -46 -191 -42
rect -207 -48 -187 -46
rect -347 -66 -342 -50
rect -343 -70 -342 -66
rect -340 -54 -338 -50
rect -334 -54 -332 -50
rect -340 -70 -332 -54
rect -330 -66 -325 -50
rect -253 -53 -237 -49
rect -253 -54 -233 -53
rect -207 -51 -187 -50
rect -203 -55 -187 -51
rect -253 -58 -233 -56
rect -249 -62 -233 -58
rect -253 -64 -233 -62
rect -203 -63 -187 -59
rect -207 -64 -187 -63
rect -330 -70 -329 -66
rect -253 -67 -233 -66
rect -253 -71 -237 -67
rect -207 -67 -187 -66
rect -207 -71 -191 -67
rect 319 -70 324 -34
rect 326 -70 334 -30
rect 336 -66 341 -30
rect 336 -70 337 -66
rect -273 -94 -237 -90
rect -273 -95 -233 -94
rect -273 -105 -233 -97
rect -273 -108 -233 -107
rect -269 -112 -233 -108
rect -273 -122 -257 -118
rect -273 -123 -253 -122
rect 9 -120 14 -84
rect 13 -124 14 -120
rect 16 -124 24 -84
rect 26 -88 27 -84
rect 26 -124 31 -88
rect 52 -119 57 -103
rect 56 -123 57 -119
rect 59 -107 61 -103
rect 65 -107 67 -103
rect 59 -123 67 -107
rect 69 -119 74 -103
rect 69 -123 70 -119
rect 78 -119 83 -103
rect 82 -123 83 -119
rect 85 -107 86 -103
rect 85 -123 90 -107
rect -273 -126 -253 -125
rect -269 -130 -253 -126
rect 13 -153 14 -149
rect 9 -189 14 -153
rect 16 -189 24 -149
rect 26 -185 31 -149
rect 72 -153 73 -149
rect 68 -169 73 -153
rect 75 -165 83 -149
rect 75 -169 77 -165
rect 81 -169 83 -165
rect 85 -153 86 -149
rect 85 -169 90 -153
rect 113 -153 114 -149
rect 26 -189 27 -185
rect 41 -173 42 -169
rect 37 -189 42 -173
rect 44 -185 49 -169
rect 44 -189 45 -185
rect 109 -189 114 -153
rect 116 -189 124 -149
rect 126 -185 131 -149
rect 126 -189 127 -185
rect 141 -173 142 -169
rect 137 -189 142 -173
rect 144 -185 149 -169
rect 144 -189 145 -185
rect -52 -245 -16 -241
rect -52 -246 -12 -245
rect 68 -245 84 -241
rect 68 -246 88 -245
rect -52 -256 -12 -248
rect 68 -250 88 -248
rect 72 -254 88 -250
rect 68 -256 88 -254
rect -52 -259 -12 -258
rect -48 -263 -12 -259
rect 68 -259 88 -258
rect 68 -263 84 -259
<< ndcontact >>
rect 4 259 8 263
rect 19 259 23 263
rect 25 250 29 254
rect -12 241 -8 245
rect 19 241 23 245
rect -58 174 -54 178
rect -40 158 -36 162
rect -17 163 -13 167
rect -9 157 -5 161
rect 51 161 55 165
rect 105 161 109 165
rect 1 150 5 154
rect 10 156 14 160
rect 19 150 23 154
rect 57 153 61 157
rect 111 153 115 157
rect 267 152 271 156
rect 57 142 61 146
rect 57 134 61 138
rect 283 134 287 138
rect 145 130 149 134
rect -240 124 -236 128
rect 139 122 143 126
rect -240 116 -236 120
rect 132 112 136 116
rect -240 105 -236 109
rect -186 105 -182 109
rect 138 103 142 107
rect -246 97 -242 101
rect -192 97 -188 101
rect 292 108 296 112
rect 132 94 136 98
rect 286 99 290 103
rect 292 90 296 94
rect -240 70 -236 74
rect 165 67 169 71
rect -240 62 -236 66
rect -240 51 -236 55
rect -186 51 -182 55
rect 267 67 271 71
rect 159 59 163 63
rect -53 50 -49 54
rect -246 43 -242 47
rect -192 43 -188 47
rect 157 51 161 55
rect 283 49 287 53
rect -45 44 -41 48
rect 141 33 145 37
rect -473 3 -469 7
rect -465 9 -461 13
rect -347 1 -343 5
rect -338 7 -334 11
rect -302 6 -298 10
rect -143 6 -139 10
rect -329 1 -325 5
rect -296 -3 -292 1
rect -149 -3 -145 1
rect 279 26 283 30
rect 319 26 323 30
rect 285 18 289 22
rect -72 -4 -68 0
rect -347 -14 -343 -10
rect -302 -12 -298 -8
rect -143 -12 -139 -8
rect -64 -4 -60 0
rect -53 -4 -49 0
rect 133 8 137 12
rect 292 8 296 12
rect 337 10 341 14
rect 139 -1 143 3
rect 286 -1 290 3
rect -45 -10 -41 -6
rect 9 -13 13 -9
rect 17 -7 21 -3
rect 319 -5 323 -1
rect 133 -10 137 -6
rect 292 -10 296 -6
rect 328 -11 332 -7
rect 337 -5 341 -1
rect -295 -22 -291 -18
rect -329 -30 -325 -26
rect -289 -30 -285 -26
rect -473 -51 -469 -47
rect -465 -45 -461 -41
rect -454 -45 -450 -41
rect -446 -45 -442 -41
rect -151 -37 -147 -33
rect -293 -53 -289 -49
rect -167 -55 -163 -51
rect 9 -59 13 -55
rect -169 -63 -165 -59
rect 18 -65 22 -61
rect 27 -59 31 -55
rect -277 -71 -273 -67
rect -175 -71 -171 -67
rect 52 -67 56 -63
rect 70 -83 74 -79
rect -302 -94 -298 -90
rect -296 -103 -292 -99
rect -302 -112 -298 -108
rect -295 -122 -291 -118
rect 78 -85 82 -81
rect 86 -91 90 -87
rect -289 -130 -285 -126
rect 9 -218 13 -214
rect 18 -212 22 -208
rect 37 -211 41 -207
rect 45 -205 49 -201
rect 68 -209 72 -205
rect 86 -193 90 -189
rect 27 -218 31 -214
rect 109 -218 113 -214
rect 118 -212 122 -208
rect 137 -211 141 -207
rect 145 -205 149 -201
rect 127 -218 131 -214
rect 13 -245 17 -241
rect 44 -245 48 -241
rect 7 -254 11 -250
rect 13 -263 17 -259
rect 28 -263 32 -259
<< pdcontact >>
rect -52 259 -48 263
rect 84 259 88 263
rect -36 250 -32 254
rect -52 241 -48 245
rect 48 241 52 245
rect -58 214 -54 218
rect -49 198 -45 202
rect -40 214 -36 218
rect -17 179 -13 183
rect -9 195 -5 199
rect 1 179 5 183
rect 19 215 23 219
rect 89 161 93 165
rect 144 161 148 165
rect 73 153 77 157
rect 128 153 132 157
rect 227 152 231 156
rect 73 142 77 146
rect 243 143 247 147
rect 73 134 77 138
rect 227 134 231 138
rect 161 130 165 134
rect -224 124 -220 128
rect 177 122 181 126
rect -224 116 -220 120
rect 161 112 165 116
rect -224 105 -220 109
rect -169 105 -165 109
rect -208 97 -204 101
rect 263 108 267 112
rect -153 97 -149 101
rect 197 94 201 98
rect 227 90 231 94
rect -347 66 -343 70
rect -473 42 -469 46
rect -224 70 -220 74
rect -53 67 -49 71
rect -45 83 -41 87
rect -224 62 -220 66
rect -224 51 -220 55
rect -169 51 -165 55
rect 181 67 185 71
rect 227 67 231 71
rect 319 66 323 70
rect 197 59 201 63
rect 243 58 247 62
rect -208 43 -204 47
rect -153 43 -149 47
rect 197 51 201 55
rect 227 49 231 53
rect 328 50 332 54
rect 337 66 341 70
rect -329 30 -325 34
rect 181 42 185 46
rect 197 33 201 37
rect -465 26 -461 30
rect -72 12 -68 16
rect -64 12 -60 16
rect -53 12 -49 16
rect -45 28 -41 32
rect 9 25 13 29
rect -237 6 -233 10
rect -208 6 -204 10
rect 263 26 267 30
rect 247 18 251 22
rect 17 9 21 13
rect -473 -13 -469 -9
rect -465 -29 -461 -25
rect -454 -29 -450 -25
rect -446 -29 -442 -25
rect -273 -12 -269 -8
rect -172 -12 -168 -8
rect 162 8 166 12
rect 263 8 267 12
rect 198 -10 202 -6
rect 227 -10 231 -6
rect -257 -22 -253 -18
rect -273 -30 -269 -26
rect -207 -37 -203 -33
rect 319 -34 323 -30
rect -191 -46 -187 -42
rect -347 -70 -343 -66
rect -338 -54 -334 -50
rect -237 -53 -233 -49
rect -207 -55 -203 -51
rect -253 -62 -249 -58
rect -207 -63 -203 -59
rect -329 -70 -325 -66
rect -237 -71 -233 -67
rect -191 -71 -187 -67
rect 337 -70 341 -66
rect -237 -94 -233 -90
rect -273 -112 -269 -108
rect -257 -122 -253 -118
rect 9 -124 13 -120
rect 27 -88 31 -84
rect 52 -123 56 -119
rect 61 -107 65 -103
rect 70 -123 74 -119
rect 78 -123 82 -119
rect 86 -107 90 -103
rect -273 -130 -269 -126
rect 9 -153 13 -149
rect 68 -153 72 -149
rect 77 -169 81 -165
rect 86 -153 90 -149
rect 109 -153 113 -149
rect 27 -189 31 -185
rect 37 -173 41 -169
rect 45 -189 49 -185
rect 127 -189 131 -185
rect 137 -173 141 -169
rect 145 -189 149 -185
rect -16 -245 -12 -241
rect 84 -245 88 -241
rect 68 -254 72 -250
rect -52 -263 -48 -259
rect 84 -263 88 -259
<< polysilicon >>
rect -56 256 -52 258
rect -32 256 -12 258
rect 8 256 11 258
rect 16 256 19 258
rect 29 256 48 258
rect 88 256 91 258
rect -56 246 -52 248
rect -32 246 -12 248
rect 8 246 11 248
rect 16 246 19 248
rect 29 246 48 248
rect 88 246 91 248
rect -53 218 -51 222
rect -43 218 -41 222
rect 6 219 8 222
rect 16 219 18 222
rect -12 199 -10 203
rect -53 178 -51 198
rect -43 178 -41 198
rect -12 167 -10 179
rect -53 155 -51 158
rect -43 155 -41 158
rect 6 160 8 179
rect 16 160 18 179
rect -12 153 -10 157
rect 48 158 51 160
rect 61 158 73 160
rect 93 158 97 160
rect 101 158 105 160
rect 115 158 128 160
rect 148 158 152 160
rect 6 147 8 150
rect 16 147 18 150
rect 223 149 227 151
rect 247 149 267 151
rect 287 149 290 151
rect 45 139 51 141
rect 61 139 64 141
rect 70 139 73 141
rect 93 139 105 141
rect 223 139 227 141
rect 247 139 267 141
rect 287 139 290 141
rect 135 127 139 129
rect 149 127 161 129
rect 181 127 185 129
rect -252 121 -246 123
rect -236 121 -233 123
rect -227 121 -224 123
rect -204 121 -192 123
rect 129 109 132 111
rect 142 109 161 111
rect 201 109 204 111
rect -249 102 -246 104
rect -236 102 -224 104
rect -204 102 -200 104
rect -196 102 -192 104
rect -182 102 -169 104
rect -149 102 -145 104
rect 224 105 227 107
rect 267 105 286 107
rect 296 105 299 107
rect 129 99 132 101
rect 142 99 161 101
rect 201 99 204 101
rect 224 95 227 97
rect 267 95 286 97
rect 296 95 299 97
rect -48 87 -46 91
rect -342 70 -340 73
rect -332 70 -330 73
rect -468 46 -466 50
rect -252 67 -246 69
rect -236 67 -233 69
rect -227 67 -224 69
rect -204 67 -192 69
rect -48 54 -46 67
rect 324 70 326 74
rect 334 70 336 74
rect 155 64 159 66
rect 169 64 181 66
rect 201 64 205 66
rect 223 64 227 66
rect 247 64 267 66
rect 287 64 290 66
rect -249 48 -246 50
rect -236 48 -224 50
rect -204 48 -200 50
rect -196 48 -192 50
rect -182 48 -169 50
rect -149 48 -145 50
rect 223 54 227 56
rect 247 54 267 56
rect 287 54 290 56
rect 138 48 141 50
rect 161 48 181 50
rect 201 48 205 50
rect -67 32 -65 44
rect -48 40 -46 44
rect 138 38 141 40
rect 161 38 181 40
rect 201 38 205 40
rect -48 32 -46 36
rect -468 13 -466 26
rect -342 11 -340 30
rect -332 11 -330 30
rect 14 29 16 33
rect 324 30 326 50
rect 334 30 336 50
rect -468 -1 -466 3
rect -468 -9 -466 -5
rect -449 -9 -447 3
rect -67 9 -65 12
rect -305 3 -302 5
rect -292 3 -273 5
rect -233 3 -230 5
rect -211 3 -208 5
rect -168 3 -149 5
rect -139 3 -136 5
rect -342 -2 -340 1
rect -332 -2 -330 1
rect -67 0 -65 3
rect -48 0 -46 12
rect 243 23 247 25
rect 267 23 279 25
rect 289 23 293 25
rect -305 -7 -302 -5
rect -292 -7 -273 -5
rect -233 -7 -230 -5
rect -211 -7 -208 -5
rect -168 -7 -149 -5
rect -139 -7 -136 -5
rect -342 -10 -340 -7
rect -332 -10 -330 -7
rect -468 -41 -466 -29
rect -449 -32 -447 -29
rect 14 -3 16 9
rect 324 7 326 10
rect 334 7 336 10
rect 130 5 133 7
rect 143 5 162 7
rect 202 5 205 7
rect 224 5 227 7
rect 267 5 286 7
rect 296 5 299 7
rect 324 -1 326 2
rect 334 -1 336 2
rect -67 -16 -65 -10
rect -48 -13 -46 -10
rect 130 -5 133 -3
rect 143 -5 162 -3
rect 202 -5 205 -3
rect 224 -5 227 -3
rect 267 -5 286 -3
rect 296 -5 299 -3
rect 14 -17 16 -13
rect -299 -25 -295 -23
rect -285 -25 -273 -23
rect -253 -25 -249 -23
rect 324 -30 326 -11
rect 334 -30 336 -11
rect -449 -41 -447 -38
rect -342 -50 -340 -30
rect -332 -50 -330 -30
rect -211 -40 -207 -38
rect -187 -40 -167 -38
rect -147 -40 -144 -38
rect -468 -54 -466 -51
rect -449 -57 -447 -51
rect -211 -50 -207 -48
rect -187 -50 -167 -48
rect -147 -50 -144 -48
rect -296 -56 -293 -54
rect -273 -56 -253 -54
rect -233 -56 -229 -54
rect 14 -55 16 -52
rect 24 -55 26 -52
rect -296 -66 -293 -64
rect -273 -66 -253 -64
rect -233 -66 -229 -64
rect -211 -66 -207 -64
rect -187 -66 -175 -64
rect -165 -66 -161 -64
rect 57 -63 59 -60
rect 67 -63 69 -60
rect -342 -74 -340 -70
rect -332 -74 -330 -70
rect 14 -84 16 -65
rect 24 -84 26 -65
rect 324 -73 326 -70
rect 334 -73 336 -70
rect 83 -81 85 -77
rect -305 -97 -302 -95
rect -292 -97 -273 -95
rect -233 -97 -230 -95
rect -305 -107 -302 -105
rect -292 -107 -273 -105
rect -233 -107 -230 -105
rect -299 -125 -295 -123
rect -285 -125 -273 -123
rect -253 -125 -249 -123
rect 57 -103 59 -83
rect 67 -103 69 -83
rect 83 -103 85 -91
rect 14 -127 16 -124
rect 24 -127 26 -124
rect 57 -127 59 -123
rect 67 -127 69 -123
rect 83 -127 85 -123
rect 14 -149 16 -146
rect 24 -149 26 -146
rect 73 -149 75 -145
rect 83 -149 85 -145
rect 114 -149 116 -146
rect 124 -149 126 -146
rect 42 -169 44 -165
rect 73 -189 75 -169
rect 83 -189 85 -169
rect 142 -169 144 -165
rect 14 -208 16 -189
rect 24 -208 26 -189
rect 42 -201 44 -189
rect 114 -208 116 -189
rect 124 -208 126 -189
rect 142 -201 144 -189
rect 42 -215 44 -211
rect 73 -212 75 -209
rect 83 -212 85 -209
rect 142 -215 144 -211
rect 14 -221 16 -218
rect 24 -221 26 -218
rect 114 -221 116 -218
rect 124 -221 126 -218
rect -55 -248 -52 -246
rect -12 -248 7 -246
rect 17 -248 20 -246
rect 25 -248 28 -246
rect 48 -248 68 -246
rect 88 -248 92 -246
rect -55 -258 -52 -256
rect -12 -258 7 -256
rect 17 -258 20 -256
rect 25 -258 28 -256
rect 48 -258 68 -256
rect 88 -258 92 -256
<< polycontact >>
rect -25 258 -21 262
rect 30 258 34 262
rect -17 248 -13 252
rect 37 248 41 252
rect -51 179 -47 183
rect -41 187 -37 191
rect -10 168 -6 172
rect 8 168 12 172
rect 18 161 22 165
rect 62 160 66 164
rect 116 160 120 164
rect 100 141 104 145
rect 262 145 266 149
rect 46 135 50 139
rect 254 135 258 139
rect -251 123 -247 127
rect 150 123 154 127
rect -197 117 -193 121
rect 150 105 154 109
rect -235 98 -231 102
rect -181 98 -177 102
rect 143 95 147 99
rect 274 101 278 105
rect 281 91 285 95
rect -251 69 -247 73
rect -197 63 -193 67
rect 170 60 174 64
rect -46 55 -42 59
rect 262 60 266 64
rect -235 44 -231 48
rect -181 44 -177 48
rect 254 50 258 54
rect -65 39 -61 43
rect 162 44 166 48
rect 170 34 174 38
rect -472 14 -468 18
rect -346 12 -342 16
rect -336 19 -332 23
rect 326 31 330 35
rect 336 39 340 43
rect -453 -2 -449 2
rect -291 5 -287 9
rect -154 5 -150 9
rect -284 -5 -280 -1
rect -161 -5 -157 -1
rect 274 19 278 23
rect -46 1 -42 5
rect -472 -40 -468 -36
rect 10 -2 14 2
rect 151 1 155 5
rect 274 1 278 5
rect -71 -15 -67 -11
rect 144 -9 148 -5
rect 281 -9 285 -5
rect -284 -23 -280 -19
rect 326 -23 330 -19
rect 336 -16 340 -12
rect -346 -43 -342 -39
rect -336 -35 -332 -31
rect -180 -38 -176 -34
rect -172 -48 -168 -44
rect -447 -56 -443 -52
rect -264 -54 -260 -50
rect -272 -64 -268 -60
rect -180 -64 -176 -60
rect 10 -70 14 -66
rect 20 -77 24 -73
rect -291 -95 -287 -91
rect -284 -105 -280 -101
rect -284 -123 -280 -119
rect 53 -96 57 -92
rect 63 -88 67 -84
rect 79 -96 83 -92
rect 69 -180 73 -176
rect 79 -188 83 -184
rect 10 -207 14 -203
rect 20 -200 24 -196
rect 38 -200 42 -196
rect 110 -207 114 -203
rect 120 -200 124 -196
rect 138 -200 142 -196
rect -5 -252 -1 -248
rect 49 -252 53 -248
rect 2 -262 6 -258
rect 57 -262 61 -258
<< metal1 >>
rect -6 278 -3 287
rect -25 275 41 278
rect -62 259 -52 263
rect -25 262 -21 275
rect -62 245 -59 259
rect -17 269 20 272
rect -32 250 -21 254
rect -25 245 -21 250
rect -17 252 -13 269
rect 25 269 34 272
rect 8 259 19 263
rect 30 262 34 269
rect 12 245 15 259
rect 29 250 34 254
rect 30 245 34 250
rect 37 252 41 275
rect 88 259 98 263
rect -62 241 -52 245
rect -25 241 -12 245
rect 12 241 19 245
rect 30 241 48 245
rect -25 234 -21 241
rect 30 235 34 241
rect -284 231 -21 234
rect -347 70 -343 80
rect -473 46 -469 56
rect -479 14 -472 18
rect -465 13 -461 26
rect -362 19 -336 23
rect -485 4 -473 7
rect -455 -2 -453 2
rect -480 -13 -473 -9
rect -362 -21 -359 19
rect -329 16 -325 30
rect -366 -24 -359 -21
rect -465 -36 -461 -29
rect -454 -36 -450 -29
rect -476 -40 -472 -36
rect -465 -41 -460 -36
rect -455 -41 -450 -36
rect -480 -60 -477 -41
rect -446 -36 -442 -29
rect -446 -40 -430 -36
rect -446 -41 -442 -40
rect -473 -52 -469 -51
rect -456 -56 -447 -52
rect -443 -56 -441 -52
rect -433 -60 -430 -40
rect -362 -39 -359 -24
rect -356 12 -346 16
rect -338 12 -317 16
rect -312 13 -287 16
rect -356 7 -353 12
rect -338 11 -334 12
rect -309 6 -302 10
rect -291 9 -287 13
rect -356 -31 -353 2
rect -347 -3 -343 1
rect -329 -3 -325 1
rect -347 -6 -325 -3
rect -347 -10 -343 -6
rect -309 -8 -306 6
rect -292 -3 -287 1
rect -291 -8 -287 -3
rect -284 -1 -281 231
rect -278 225 -101 228
rect -278 27 -275 225
rect -58 225 -36 228
rect -58 218 -54 225
rect -40 218 -36 225
rect -49 191 -45 198
rect -28 191 -25 231
rect -9 226 23 229
rect -9 199 -5 226
rect 19 219 23 226
rect -60 187 -45 191
rect -37 187 -25 191
rect -60 186 -54 187
rect -64 151 -61 186
rect -58 178 -54 186
rect -47 179 -27 183
rect -30 172 -27 179
rect -17 172 -13 179
rect 1 172 5 179
rect 30 172 34 230
rect -30 168 -13 172
rect -6 168 5 172
rect 12 168 34 172
rect 39 169 61 172
rect -17 167 -13 168
rect 1 165 5 168
rect 1 161 14 165
rect 22 161 31 165
rect -40 155 -36 158
rect -64 148 -12 151
rect -258 137 -231 140
rect -258 93 -255 137
rect -251 127 -247 129
rect -235 128 -231 137
rect -236 124 -224 128
rect -251 114 -247 123
rect -236 116 -224 120
rect -236 115 -231 116
rect -197 115 -193 117
rect -236 109 -231 110
rect -236 105 -224 109
rect -182 105 -169 109
rect -247 97 -246 101
rect -235 94 -231 98
rect -258 90 -236 93
rect -208 90 -204 97
rect -208 87 -198 90
rect -258 83 -231 86
rect -191 85 -188 97
rect -181 91 -177 98
rect -149 97 -139 101
rect -45 87 -41 97
rect -258 39 -255 83
rect -251 73 -247 75
rect -235 74 -231 83
rect -236 70 -224 74
rect -251 60 -247 69
rect -236 62 -224 66
rect -236 61 -231 62
rect -197 61 -193 63
rect -236 55 -231 56
rect -236 51 -224 55
rect -182 51 -169 55
rect -53 54 -49 67
rect -42 55 -35 59
rect -247 43 -246 47
rect -235 40 -231 44
rect -258 36 -236 39
rect -208 36 -204 43
rect -208 33 -198 36
rect -191 31 -188 43
rect -181 37 -177 44
rect -149 43 -139 47
rect -34 45 -31 54
rect -61 39 -59 43
rect -45 39 -41 44
rect -34 32 -31 40
rect -41 28 -31 32
rect -278 24 -150 27
rect -233 6 -223 10
rect -218 6 -208 10
rect -309 -12 -302 -8
rect -291 -12 -273 -8
rect -309 -18 -306 -12
rect -309 -22 -295 -18
rect -284 -19 -280 -12
rect -226 -18 -223 6
rect -161 -1 -157 16
rect -153 13 -150 24
rect -154 9 -150 13
rect -139 6 -132 10
rect -154 -3 -149 1
rect -154 -8 -150 -3
rect -135 -8 -132 6
rect -72 5 -68 12
rect -168 -12 -150 -8
rect -139 -12 -132 -8
rect -84 1 -68 5
rect -253 -22 -223 -18
rect -154 -19 -150 -12
rect -180 -22 -150 -19
rect -84 -19 -81 1
rect -72 0 -68 1
rect -64 5 -60 12
rect -53 5 -49 12
rect -64 0 -59 5
rect -54 0 -49 5
rect -42 1 -38 5
rect -45 -11 -41 -10
rect -73 -15 -71 -11
rect -67 -15 -58 -11
rect -37 -19 -34 0
rect -15 -12 -12 148
rect -9 146 -5 157
rect 10 160 14 161
rect 1 146 5 150
rect 19 146 23 150
rect -9 143 23 146
rect 28 49 31 161
rect 39 125 42 169
rect 50 161 51 165
rect 62 164 66 168
rect 89 172 101 175
rect 89 165 93 172
rect 106 172 115 175
rect 100 161 105 165
rect 116 164 120 171
rect 148 161 158 165
rect 61 153 73 157
rect 115 153 128 157
rect 254 156 258 162
rect 46 139 50 148
rect 61 152 66 153
rect 61 146 66 147
rect 217 152 227 156
rect 254 152 267 156
rect 61 142 73 146
rect 100 145 104 147
rect 150 141 211 144
rect 46 133 50 135
rect 61 134 73 138
rect 150 134 154 141
rect 62 125 66 134
rect 149 130 161 134
rect 208 132 211 141
rect 217 138 220 152
rect 254 147 258 152
rect 247 143 258 147
rect 217 135 227 138
rect 208 129 217 132
rect 214 127 217 129
rect 254 127 258 135
rect 39 122 66 125
rect 125 122 139 126
rect 125 116 128 122
rect 150 116 154 123
rect 181 122 211 126
rect 214 124 258 127
rect 125 112 132 116
rect 143 112 161 116
rect 125 98 128 112
rect 143 107 147 112
rect 142 103 147 107
rect 125 94 132 98
rect 143 69 147 95
rect 150 88 154 105
rect 208 98 211 122
rect 262 123 266 145
rect 287 134 290 138
rect 262 120 278 123
rect 274 112 278 120
rect 267 108 285 112
rect 296 108 303 112
rect 201 94 211 98
rect 217 90 227 94
rect 274 83 278 101
rect 281 103 285 108
rect 281 99 286 103
rect 170 80 278 83
rect 300 94 303 108
rect 170 71 174 80
rect 281 77 285 91
rect 296 90 303 94
rect 259 74 285 77
rect 319 77 341 80
rect 254 71 259 72
rect 128 66 147 69
rect 169 67 181 71
rect 217 67 227 71
rect 254 67 267 71
rect 319 70 323 77
rect 128 49 131 66
rect 28 46 131 49
rect 134 59 159 63
rect 9 29 13 39
rect 17 2 21 9
rect 28 2 31 46
rect 134 37 137 59
rect 170 55 174 60
rect 201 59 211 63
rect 208 55 211 59
rect 161 51 174 55
rect 201 51 211 55
rect 134 33 141 37
rect 162 28 166 44
rect 170 46 174 51
rect 170 42 181 46
rect 131 25 166 28
rect 208 37 211 51
rect 217 53 220 67
rect 254 62 258 67
rect 337 70 341 77
rect 247 58 258 62
rect 217 49 227 53
rect 254 40 258 50
rect 262 46 266 60
rect 287 49 290 53
rect 262 43 284 46
rect 281 40 307 43
rect 254 37 278 40
rect 328 43 332 50
rect 312 39 332 43
rect 340 39 356 43
rect 170 22 174 34
rect 201 33 211 37
rect 274 30 278 37
rect 319 30 323 39
rect 330 31 350 35
rect 267 26 279 30
rect 144 19 174 22
rect 144 12 148 19
rect 217 18 247 22
rect -2 -2 10 2
rect 17 -2 31 2
rect 126 8 133 12
rect 144 8 162 12
rect -84 -22 -34 -19
rect -285 -30 -273 -26
rect -356 -35 -336 -31
rect -329 -39 -325 -30
rect -284 -37 -280 -30
rect -217 -37 -207 -33
rect -180 -34 -176 -22
rect -2 -25 1 -2
rect 17 -3 21 -2
rect 126 -6 129 8
rect 144 3 148 8
rect 143 -1 148 3
rect 126 -10 133 -6
rect 9 -17 13 -13
rect 144 -13 148 -9
rect 144 -25 147 -13
rect 151 -16 155 1
rect 217 -6 220 18
rect 274 12 278 19
rect 289 18 303 22
rect 300 12 303 18
rect 267 8 285 12
rect 296 8 303 12
rect 202 -10 212 -6
rect 217 -10 227 -6
rect -362 -43 -346 -39
rect -338 -43 -318 -39
rect -338 -50 -334 -43
rect -284 -40 -260 -37
rect -313 -43 -287 -40
rect -290 -46 -268 -43
rect -296 -53 -293 -49
rect -480 -63 -430 -60
rect -272 -60 -268 -46
rect -264 -50 -260 -40
rect -233 -53 -223 -49
rect -264 -62 -253 -58
rect -347 -77 -343 -70
rect -264 -67 -260 -62
rect -226 -67 -223 -53
rect -217 -51 -214 -37
rect -172 -28 1 -25
rect -187 -46 -176 -42
rect -180 -51 -176 -46
rect -172 -44 -168 -28
rect -147 -37 -140 -33
rect -217 -55 -207 -51
rect -180 -55 -167 -51
rect -217 -59 -214 -55
rect -217 -63 -207 -59
rect -180 -60 -176 -55
rect -143 -59 -140 -37
rect 9 -51 31 -48
rect 9 -55 13 -51
rect 27 -55 31 -51
rect -165 -63 -140 -59
rect 18 -66 22 -65
rect -329 -77 -325 -70
rect -273 -70 -260 -67
rect -273 -71 -268 -70
rect -347 -80 -325 -77
rect -291 -75 -268 -74
rect -263 -75 -260 -70
rect -233 -71 -223 -67
rect -187 -71 -175 -67
rect -9 -69 10 -66
rect -291 -77 -260 -75
rect -309 -94 -302 -90
rect -291 -91 -287 -77
rect -180 -80 -176 -71
rect -9 -77 -6 -69
rect 6 -70 10 -69
rect 18 -70 41 -66
rect 3 -77 20 -73
rect -309 -108 -306 -94
rect -284 -83 -176 -80
rect -292 -103 -287 -99
rect -291 -108 -287 -103
rect -284 -101 -280 -83
rect 27 -84 31 -70
rect -233 -94 -223 -90
rect -309 -112 -302 -108
rect -291 -112 -273 -108
rect -309 -118 -306 -112
rect -309 -122 -295 -118
rect -284 -119 -280 -112
rect -226 -118 -223 -94
rect 38 -92 41 -70
rect 44 -84 47 -52
rect 52 -59 82 -56
rect 52 -63 56 -59
rect 44 -88 63 -84
rect 70 -92 74 -83
rect 78 -81 82 -59
rect 86 -92 90 -91
rect 38 -96 53 -92
rect 61 -96 79 -92
rect 86 -96 102 -92
rect 61 -103 65 -96
rect 86 -103 90 -96
rect -253 -122 -223 -118
rect -285 -130 -273 -126
rect -284 -136 -280 -130
rect 9 -134 13 -124
rect 52 -130 56 -123
rect 70 -130 74 -123
rect 78 -130 82 -123
rect 52 -133 82 -130
rect 9 -142 41 -139
rect 9 -149 13 -142
rect 37 -169 41 -142
rect 68 -142 90 -139
rect 68 -149 72 -142
rect 86 -149 90 -142
rect 77 -176 81 -169
rect 56 -180 69 -176
rect 77 -180 96 -176
rect 27 -196 31 -189
rect 45 -196 49 -189
rect 56 -196 59 -180
rect -311 -200 20 -197
rect 27 -200 38 -196
rect 45 -200 59 -196
rect 62 -188 79 -184
rect 27 -203 31 -200
rect 3 -207 10 -203
rect 18 -207 31 -203
rect 45 -201 49 -200
rect 62 -203 65 -188
rect 86 -189 90 -180
rect 59 -206 65 -203
rect 93 -203 96 -180
rect 99 -196 102 -96
rect 109 -142 141 -139
rect 109 -149 113 -142
rect 137 -169 141 -142
rect 127 -196 131 -189
rect 145 -196 149 -189
rect 99 -200 120 -196
rect 127 -200 138 -196
rect 145 -200 155 -196
rect 127 -203 131 -200
rect 3 -228 6 -207
rect 18 -208 22 -207
rect 9 -222 13 -218
rect 27 -222 31 -218
rect 37 -222 41 -211
rect 9 -225 41 -222
rect 59 -226 62 -206
rect 93 -207 110 -203
rect 118 -207 131 -203
rect 145 -201 149 -200
rect 68 -212 72 -209
rect 118 -208 122 -207
rect 109 -222 113 -218
rect 127 -222 131 -218
rect 137 -222 141 -211
rect 109 -225 141 -222
rect 58 -228 62 -226
rect 275 -228 278 1
rect 281 3 285 8
rect 281 -1 286 3
rect 300 -6 303 8
rect 337 6 341 10
rect 319 3 341 6
rect 319 -1 323 3
rect 337 -1 341 3
rect 347 -2 350 31
rect 281 -13 285 -9
rect 296 -10 303 -6
rect 328 -12 332 -11
rect 347 -12 350 -7
rect 281 -16 306 -13
rect 311 -16 332 -12
rect 340 -16 350 -12
rect 353 24 356 39
rect 353 21 365 24
rect 319 -30 323 -16
rect 353 -19 356 21
rect 330 -23 356 -19
rect 337 -80 341 -70
rect 58 -231 278 -228
rect 2 -241 6 -233
rect 58 -235 61 -231
rect 57 -241 61 -235
rect -12 -245 6 -241
rect 17 -245 24 -241
rect 48 -245 61 -241
rect 88 -245 98 -241
rect -62 -263 -52 -259
rect -5 -275 -1 -252
rect 2 -250 6 -245
rect 2 -254 7 -250
rect 21 -259 24 -245
rect 2 -269 6 -262
rect 17 -263 28 -259
rect 2 -272 11 -269
rect 49 -269 53 -252
rect 57 -250 61 -245
rect 57 -254 68 -250
rect 16 -272 53 -269
rect 95 -259 98 -245
rect 57 -275 61 -262
rect 88 -263 98 -259
rect -5 -278 61 -275
rect 39 -287 42 -278
<< m2contact >>
rect 20 267 25 272
rect -484 13 -479 18
rect -461 14 -456 19
rect -485 -14 -480 -9
rect -474 -57 -469 -52
rect -461 -57 -456 -52
rect -441 -57 -436 -52
rect -317 12 -312 17
rect -356 2 -351 7
rect -101 223 -96 228
rect 29 230 34 235
rect -65 186 -60 191
rect -252 129 -247 134
rect -252 109 -247 114
rect -181 109 -176 114
rect -252 96 -247 101
rect -182 86 -177 91
rect -252 75 -247 80
rect -252 55 -247 60
rect -181 55 -176 60
rect -58 55 -53 60
rect -35 54 -30 59
rect -252 42 -247 47
rect -182 32 -177 37
rect -161 16 -156 21
rect -78 -16 -73 -11
rect -58 -16 -53 -11
rect -45 -16 -40 -11
rect 45 161 50 166
rect 115 171 120 176
rect 45 148 50 153
rect 116 148 121 153
rect 45 128 50 133
rect 254 72 259 77
rect 126 25 131 30
rect 307 39 312 44
rect -16 -17 -11 -12
rect 150 -21 155 -16
rect -318 -44 -313 -39
rect 142 -30 147 -25
rect 43 -52 48 -47
rect -268 -75 -263 -70
rect -2 -77 3 -72
rect -11 -82 -6 -77
rect -316 -200 -311 -195
rect 345 -7 350 -2
rect 306 -17 311 -12
rect 2 -233 7 -228
rect 11 -272 16 -267
<< metal2 >>
rect 21 272 24 287
rect -99 230 29 233
rect -99 228 -96 230
rect -172 186 -65 189
rect -247 130 -177 133
rect -180 114 -177 130
rect -251 101 -247 109
rect -198 87 -197 90
rect -192 87 -182 90
rect -172 89 -169 186
rect 46 153 50 161
rect 117 132 120 148
rect 50 129 120 132
rect -177 86 -169 89
rect 150 81 154 88
rect -247 76 -177 79
rect 150 78 259 81
rect -180 60 -177 76
rect 254 77 259 78
rect -77 56 -58 59
rect -251 47 -247 55
rect -198 33 -197 36
rect -192 33 -182 36
rect -180 28 -177 32
rect -371 25 -177 28
rect -456 15 -437 18
rect -483 3 -480 13
rect -483 -9 -480 -2
rect -440 -52 -437 15
rect -371 6 -368 25
rect -316 17 -161 20
rect -317 9 -306 12
rect -371 3 -356 6
rect -469 -56 -461 -52
rect -316 -195 -313 -44
rect -309 -79 -306 9
rect -77 -11 -74 56
rect -23 40 129 43
rect -53 -15 -45 -11
rect -23 -72 -20 40
rect 126 30 129 40
rect 350 -6 365 -3
rect -15 -31 -12 -17
rect 155 -20 310 -17
rect 147 -28 275 -25
rect -15 -34 47 -31
rect 44 -47 47 -34
rect -263 -75 -20 -72
rect -309 -82 -11 -79
rect -1 -232 2 -77
rect 272 -230 275 -28
rect 7 -233 275 -230
rect 12 -287 15 -272
<< m3contact >>
rect -197 87 -192 92
rect -197 33 -192 38
rect -483 -2 -478 3
<< m123contact >>
rect -236 110 -231 115
rect -197 110 -192 115
rect -236 89 -231 94
rect 61 168 66 173
rect 101 170 106 175
rect 61 147 66 152
rect 100 147 105 152
rect -236 56 -231 61
rect -197 56 -192 61
rect -236 35 -231 40
rect -460 -2 -455 3
rect -481 -41 -476 -36
rect -460 -41 -455 -36
rect -371 -25 -366 -20
rect -59 39 -54 44
rect -36 40 -31 45
rect -59 0 -54 5
rect -38 0 -33 5
<< metal3 >>
rect 63 173 66 176
rect 101 152 105 170
rect -234 115 -231 144
rect 63 119 66 147
rect -196 92 -193 110
rect -234 61 -231 89
rect -196 38 -193 56
rect -54 40 -36 44
rect -234 25 -231 35
rect -369 22 -231 25
rect -478 -1 -460 2
rect -369 -20 -366 22
rect -87 2 -59 5
rect -33 2 -30 5
rect -484 -39 -481 -36
rect -455 -39 -427 -36
<< labels >>
rlabel metal1 -1 -1 1 1 1 C0
rlabel metal1 4 -1 6 1 3 in
rlabel metal1 10 -16 12 -14 1 gnd
rlabel metal1 10 36 12 38 5 vdd
rlabel metal1 24 -1 26 1 1 C0_bar
rlabel metal1 -22 169 -20 171 3 out
rlabel metal1 25 162 26 163 7 a
rlabel metal1 23 169 25 171 7 b
rlabel metal1 21 226 22 228 5 vdd
rlabel metal1 12 144 13 145 1 gnd
rlabel metal1 -24 237 -22 239 1 G0_bar
rlabel metal1 31 237 33 239 1 P0_bar
rlabel metal1 -5 279 -4 282 1 A0
rlabel metal2 22 279 23 282 1 B0
rlabel metal1 9 260 10 262 7 gnd
rlabel metal1 -61 251 -60 253 3 vdd
rlabel metal1 13 252 14 253 3 gnd
rlabel metal1 95 261 97 262 7 vdd
rlabel metal1 -337 -79 -335 -78 1 vdd
rlabel metal1 -337 -5 -336 -4 1 gnd
rlabel metal1 -346 77 -345 79 5 vdd
rlabel metal1 -346 -9 -344 -8 5 gnd
rlabel metal2 -366 4 -363 5 1 B1
rlabel metal1 -366 -23 -363 -22 1 A1
rlabel metal1 -323 13 -321 15 1 P1_bar
rlabel metal1 -323 -42 -321 -40 1 G1_bar
rlabel metal1 -34 189 -32 190 7 a
rlabel metal1 -35 180 -34 182 7 b
rlabel metal1 -39 156 -37 157 1 gnd
rlabel m2contact -62 188 -60 190 3 C1
rlabel metal1 -48 226 -46 227 5 vdd
rlabel metal1 26 -262 27 -260 3 gnd
rlabel metal1 96 -253 97 -251 7 vdd
rlabel metal1 22 -253 23 -252 7 gnd
rlabel metal1 -61 -262 -59 -261 3 vdd
rlabel metal2 13 -282 14 -282 1 B2
rlabel metal1 40 -282 41 -279 1 A2
rlabel metal1 58 -239 60 -237 1 G2_bar
rlabel metal1 3 -239 5 -237 1 P2_bar
rlabel metal1 119 -224 120 -223 1 gnd
rlabel metal1 110 -142 111 -140 5 vdd
rlabel metal1 107 -199 109 -197 3 b
rlabel metal1 106 -206 107 -205 3 a
rlabel metal1 93 -95 95 -93 7 out
rlabel metal1 53 -62 55 -61 5 gnd
rlabel metal1 50 -87 51 -85 3 b
rlabel metal1 48 -95 50 -94 3 a
rlabel metal1 62 -132 64 -131 1 vdd
rlabel metal1 19 -50 20 -49 5 gnd
rlabel metal1 10 -133 11 -131 1 vdd
rlabel metal1 33 -69 35 -67 7 out
rlabel metal1 7 -76 9 -74 3 b
rlabel metal1 6 -68 7 -67 3 a
rlabel metal1 69 -211 71 -210 1 gnd
rlabel metal1 92 -179 94 -177 1 out
rlabel metal1 66 -187 67 -185 3 b
rlabel metal1 64 -178 66 -177 3 a
rlabel metal1 78 -141 80 -140 5 vdd
rlabel metal1 52 -199 54 -197 7 out
rlabel metal1 6 -206 7 -205 3 a
rlabel metal1 7 -199 9 -197 3 b
rlabel metal1 10 -142 11 -140 5 vdd
rlabel metal1 19 -224 20 -223 1 gnd
rlabel pdiffusion 20 -178 22 -160 1 P2_bar--OR--G1_bar
rlabel pdiffusion 19 -109 22 -99 1 P2_bar--NOR--P1_bar
rlabel pdiffusion 63 -117 66 -110 1 node24--AND--C1
rlabel pdiffusion 78 -162 80 -156 1 G2_bar--AND--node24
rlabel pdiffusion 120 -174 122 -163 1 node25--OR--node23
rlabel metal1 357 22 360 23 5 A1
rlabel metal2 357 -5 360 -4 5 B1
rlabel metal1 338 8 340 9 1 gnd
rlabel metal1 339 -79 340 -77 1 vdd
rlabel metal1 330 4 331 5 5 gnd
rlabel metal1 329 78 331 79 5 vdd
rlabel metal1 -307 -1 -306 0 3 gnd
rlabel pdiffusion -258 -103 -247 -101 1 node15--OR--node13
rlabel metal1 -283 -135 -281 -133 1 C2
rlabel metal1 -308 -101 -307 -100 3 gnd
rlabel metal1 -226 -92 -224 -91 7 vdd
rlabel metal1 -283 -90 -281 -88 5 b
rlabel metal1 -290 -88 -289 -87 5 a
rlabel pdiffusion -246 -61 -240 -59 1 G1_bar--NAND--node12
rlabel pdiffusion -201 -47 -194 -44 1 node14--AND--C0
rlabel pdiffusion -193 -3 -183 0 1 P1_bar--NOR--P0_bar
rlabel pdiffusion -262 -3 -244 -1 1 P1_bar--OR--G0_bar
rlabel metal1 -179 -76 -177 -74 1 out
rlabel metal1 -146 -36 -145 -34 7 gnd
rlabel metal1 -171 -32 -169 -31 5 b
rlabel metal1 -179 -31 -178 -29 5 a
rlabel metal1 -216 -45 -215 -43 3 vdd
rlabel metal1 -134 -1 -133 0 7 gnd
rlabel metal1 -217 8 -215 9 3 vdd
rlabel metal1 -153 -16 -151 -14 1 out
rlabel metal1 -160 10 -158 12 5 b
rlabel metal1 -152 12 -151 13 5 a
rlabel metal1 -295 -52 -294 -50 3 gnd
rlabel metal1 -263 -75 -261 -73 3 out
rlabel metal1 -271 -48 -269 -47 5 b
rlabel metal1 -262 -47 -261 -45 5 a
rlabel metal1 -225 -61 -224 -59 7 vdd
rlabel metal1 -283 -35 -281 -33 1 out
rlabel metal1 -290 12 -289 13 5 a
rlabel metal1 -283 10 -281 12 5 b
rlabel metal1 -226 8 -224 9 7 vdd
rlabel metal1 301 100 302 101 7 gnd
rlabel metal1 218 91 220 92 3 vdd
rlabel metal1 275 88 277 90 1 b
rlabel metal1 283 87 284 88 1 a
rlabel metal1 171 74 173 76 5 out
rlabel metal1 139 34 140 36 3 gnd
rlabel metal1 163 31 165 32 1 b
rlabel metal1 172 29 173 31 1 a
rlabel metal1 209 43 210 45 7 vdd
rlabel metal1 127 0 128 1 3 gnd
rlabel metal1 209 -9 211 -8 7 vdd
rlabel metal1 145 14 147 16 5 out
rlabel metal1 152 -12 154 -10 1 b
rlabel metal1 145 -13 146 -12 1 a
rlabel metal1 288 50 289 52 7 gnd
rlabel metal1 263 47 265 48 1 b
rlabel metal1 255 45 256 47 1 a
rlabel metal1 218 59 219 61 3 vdd
rlabel metal1 275 33 277 35 5 out
rlabel metal1 283 -13 284 -12 1 a
rlabel metal1 275 -12 277 -10 1 b
rlabel metal1 218 -9 220 -8 3 vdd
rlabel metal1 315 -15 317 -13 1 P3_bar
rlabel metal1 315 40 317 42 1 G3_bar
rlabel pdiffusion 238 1 256 3 1 P3_bar--OR--G2_bar
rlabel pdiffusion 177 0 187 3 1 P3_bar--NOR--P2_bar
rlabel pdiffusion 188 44 195 47 1 node34--AND--node13
rlabel pdiffusion 234 59 240 61 1 node34--NAND--node14
rlabel pdiffusion 241 101 252 103 1 node33--NOR--node35
rlabel metal1 152 -199 154 -197 1 C3
rlabel m2contact 255 73 257 75 1 Pout_bar
rlabel metal1 275 114 277 117 1 Gout_bar
rlabel metal1 144 91 145 92 1 a
rlabel metal1 151 92 153 94 1 b
rlabel metal1 208 95 210 96 7 vdd
rlabel metal1 126 104 127 105 3 gnd
rlabel metal1 151 137 153 139 1 node36
rlabel metal1 218 144 219 146 3 vdd
rlabel metal1 255 130 256 132 1 a
rlabel metal1 263 132 265 133 1 b
rlabel metal1 288 135 289 137 7 gnd
rlabel metal1 255 158 257 160 1 Cout
rlabel metal1 -234 38 -232 40 3 b
rlabel metal1 -234 56 -232 60 3 out
rlabel metal1 -478 15 -476 17 3 a
rlabel metal1 -478 -39 -476 -37 1 b
rlabel metal1 -472 53 -470 55 5 vdd
rlabel metal1 -460 -39 -456 -37 1 out
rlabel metal1 -464 15 -462 18 1 a_bar
rlabel metal1 -234 92 -232 94 3 b
rlabel metal3 -233 141 -232 143 1 S1
rlabel metal1 -38 56 -36 58 7 a
rlabel metal1 -38 2 -36 4 1 b
rlabel metal1 -44 39 -42 40 1 gnd
rlabel metal1 -44 94 -42 96 5 vdd
rlabel metal1 -58 2 -54 4 1 out
rlabel metal1 -52 56 -50 59 1 a_bar
rlabel metal1 117 168 119 170 5 a
rlabel metal1 63 168 65 170 3 b
rlabel metal1 100 162 101 164 3 gnd
rlabel metal1 155 162 157 164 7 vdd
rlabel metal1 63 148 65 152 3 out
rlabel metal1 117 154 120 156 3 a_bar
rlabel metal1 -478 5 -476 6 1 gnd
rlabel metal1 -190 38 -189 40 3 gnd
rlabel metal1 -180 52 -177 54 3 a_bar
rlabel metal1 -142 44 -140 46 7 vdd
rlabel metal1 -180 38 -178 40 1 a
rlabel metal1 -190 92 -189 94 3 gnd
rlabel metal1 -180 106 -177 108 3 a_bar
rlabel metal1 -142 98 -140 100 7 vdd
rlabel metal1 -180 92 -178 94 1 a
<< end >>
