magic
tech scmos
timestamp 1731437957
<< nwell >>
rect -58 235 -26 269
rect 42 235 94 269
rect -64 192 -30 224
rect -23 173 29 225
rect 70 151 94 183
rect -199 106 -167 130
rect -144 106 -112 149
rect 51 96 94 128
rect -353 24 -319 76
rect -199 41 -167 65
rect -144 41 -112 84
rect -57 63 -33 95
rect 155 88 207 140
rect 221 128 253 162
rect 221 84 273 119
rect -279 -36 -227 16
rect -214 -18 -162 16
rect -76 8 -33 40
rect 3 3 27 35
rect 175 27 207 77
rect 221 43 253 77
rect 313 44 347 76
rect 45 -9 77 25
rect 156 -16 208 18
rect 221 -16 273 36
rect -353 -76 -319 -44
rect -259 -77 -227 -43
rect -213 -77 -181 -27
rect 94 -75 137 -43
rect 313 -76 347 -24
rect -279 -136 -227 -84
rect -190 -135 -158 -92
rect -135 -140 -103 -92
rect -80 -140 -48 -97
rect 3 -130 37 -78
rect 46 -129 96 -97
rect 113 -130 137 -98
rect 170 -142 194 -110
rect 3 -195 55 -143
rect 62 -175 96 -143
rect 103 -195 155 -143
rect 170 -197 213 -165
rect -58 -269 -6 -235
rect 62 -269 94 -235
<< ntransistor >>
rect -12 256 8 258
rect 19 256 29 258
rect -12 246 8 248
rect 19 246 29 248
rect -53 158 -51 178
rect -43 158 -41 178
rect -12 157 -10 167
rect 6 150 8 160
rect 16 150 18 160
rect 267 149 287 151
rect -106 136 -96 138
rect 81 134 83 144
rect 267 139 287 141
rect 139 127 149 129
rect -160 117 -150 119
rect -106 117 -96 119
rect 132 109 142 111
rect 286 105 296 107
rect 132 99 142 101
rect 286 95 296 97
rect -106 71 -96 73
rect 62 80 64 90
rect 81 80 83 90
rect 159 64 169 66
rect 267 64 287 66
rect -160 52 -150 54
rect -106 52 -96 54
rect -46 46 -44 56
rect 267 54 287 56
rect 141 48 161 50
rect 141 38 161 40
rect -342 1 -340 11
rect -332 1 -330 11
rect -302 3 -292 5
rect -149 3 -139 5
rect 279 23 289 25
rect 91 12 111 14
rect -302 -7 -292 -5
rect -149 -7 -139 -5
rect -342 -30 -340 -10
rect -332 -30 -330 -10
rect -65 -8 -63 2
rect -46 -8 -44 2
rect 324 10 326 30
rect 334 10 336 30
rect 133 5 143 7
rect 286 5 296 7
rect 91 2 111 4
rect 14 -13 16 -3
rect 133 -5 143 -3
rect 286 -5 296 -3
rect 324 -11 326 -1
rect 334 -11 336 -1
rect -295 -25 -285 -23
rect 105 -37 107 -27
rect 124 -37 126 -27
rect -167 -40 -147 -38
rect -167 -50 -147 -48
rect -293 -56 -273 -54
rect -293 -66 -273 -64
rect -175 -66 -165 -64
rect 14 -65 16 -55
rect 24 -65 26 -55
rect 57 -83 59 -63
rect 67 -83 69 -63
rect -302 -97 -292 -95
rect -206 -105 -196 -103
rect -152 -105 -142 -103
rect -302 -107 -292 -105
rect -42 -110 -32 -108
rect -295 -125 -285 -123
rect -206 -124 -196 -122
rect 83 -91 85 -81
rect 124 -91 126 -81
rect -96 -129 -86 -127
rect -42 -129 -32 -127
rect 181 -159 183 -149
rect 14 -218 16 -208
rect 24 -218 26 -208
rect 42 -211 44 -201
rect 73 -209 75 -189
rect 83 -209 85 -189
rect 114 -218 116 -208
rect 124 -218 126 -208
rect 142 -211 144 -201
rect 181 -213 183 -203
rect 200 -213 202 -203
rect 7 -248 17 -246
rect 28 -248 48 -246
rect 7 -258 17 -256
rect 28 -258 48 -256
<< ptransistor >>
rect -52 256 -32 258
rect 48 256 88 258
rect -52 246 -32 248
rect 48 246 88 248
rect -53 198 -51 218
rect -43 198 -41 218
rect -12 179 -10 199
rect 6 179 8 219
rect 16 179 18 219
rect 81 157 83 177
rect 227 149 247 151
rect -138 136 -118 138
rect 227 139 247 141
rect 161 127 181 129
rect -193 117 -173 119
rect -138 117 -118 119
rect 62 102 64 122
rect 81 102 83 122
rect 161 109 201 111
rect 227 105 267 107
rect 161 99 201 101
rect 227 95 267 97
rect -138 71 -118 73
rect -342 30 -340 70
rect -332 30 -330 70
rect -46 69 -44 89
rect 181 64 201 66
rect 227 64 247 66
rect -193 52 -173 54
rect -138 52 -118 54
rect 227 54 247 56
rect 181 48 201 50
rect 324 50 326 70
rect 334 50 336 70
rect 181 38 201 40
rect -65 14 -63 34
rect -46 14 -44 34
rect -273 3 -233 5
rect -208 3 -168 5
rect 14 9 16 29
rect 247 23 267 25
rect 51 12 71 14
rect -273 -7 -233 -5
rect -208 -7 -168 -5
rect 162 5 202 7
rect 227 5 267 7
rect 51 2 71 4
rect 162 -5 202 -3
rect 227 -5 267 -3
rect -273 -25 -253 -23
rect -207 -40 -187 -38
rect -342 -70 -340 -50
rect -332 -70 -330 -50
rect -207 -50 -187 -48
rect -253 -56 -233 -54
rect -253 -66 -233 -64
rect -207 -66 -187 -64
rect 105 -69 107 -49
rect 124 -69 126 -49
rect 324 -70 326 -30
rect 334 -70 336 -30
rect -273 -97 -233 -95
rect -184 -105 -164 -103
rect -129 -105 -109 -103
rect -273 -107 -233 -105
rect -74 -110 -54 -108
rect -273 -125 -253 -123
rect -184 -124 -164 -122
rect 14 -124 16 -84
rect 24 -124 26 -84
rect 57 -123 59 -103
rect 67 -123 69 -103
rect 83 -123 85 -103
rect 124 -124 126 -104
rect -129 -129 -109 -127
rect -74 -129 -54 -127
rect 181 -136 183 -116
rect 14 -189 16 -149
rect 24 -189 26 -149
rect 73 -169 75 -149
rect 83 -169 85 -149
rect 42 -189 44 -169
rect 114 -189 116 -149
rect 124 -189 126 -149
rect 142 -189 144 -169
rect 181 -191 183 -171
rect 200 -191 202 -171
rect -52 -248 -12 -246
rect 68 -248 88 -246
rect -52 -258 -12 -256
rect 68 -258 88 -256
<< ndiffusion >>
rect -12 259 4 263
rect -12 258 8 259
rect 23 259 29 263
rect 19 258 29 259
rect -12 248 8 256
rect 19 254 29 256
rect 19 250 25 254
rect 19 248 29 250
rect -12 245 8 246
rect -8 241 8 245
rect 19 245 29 246
rect 23 241 29 245
rect -54 174 -53 178
rect -58 158 -53 174
rect -51 158 -43 178
rect -41 162 -36 178
rect -41 158 -40 162
rect -13 163 -12 167
rect -17 157 -12 163
rect -10 161 -5 167
rect -10 157 -9 161
rect 1 154 6 160
rect 5 150 6 154
rect 8 156 10 160
rect 14 156 16 160
rect 8 150 16 156
rect 18 154 23 160
rect 18 150 19 154
rect 271 152 287 156
rect 267 151 287 152
rect -102 139 -96 143
rect -106 138 -96 139
rect 80 140 81 144
rect -106 135 -96 136
rect -102 131 -96 135
rect 76 134 81 140
rect 83 138 88 144
rect 267 141 287 149
rect 83 134 84 138
rect 267 138 287 139
rect 267 134 283 138
rect -156 120 -150 124
rect -160 119 -150 120
rect -102 120 -96 124
rect 139 130 145 134
rect 139 129 149 130
rect 139 126 149 127
rect 143 122 149 126
rect -106 119 -96 120
rect -160 116 -150 117
rect -160 112 -154 116
rect -106 116 -96 117
rect -106 112 -100 116
rect 136 112 142 116
rect 132 111 142 112
rect 132 107 142 109
rect 132 103 138 107
rect 132 101 142 103
rect 286 108 292 112
rect 286 107 296 108
rect 132 98 142 99
rect 136 94 142 98
rect 286 103 296 105
rect 290 99 296 103
rect 286 97 296 99
rect 286 94 296 95
rect 286 90 292 94
rect -102 74 -96 78
rect -106 73 -96 74
rect -106 70 -96 71
rect -102 66 -96 70
rect 61 86 62 90
rect 57 80 62 86
rect 64 86 65 90
rect 64 80 69 86
rect 80 86 81 90
rect 76 80 81 86
rect 83 84 88 90
rect 83 80 84 84
rect -156 55 -150 59
rect -160 54 -150 55
rect -102 55 -96 59
rect 159 67 165 71
rect 159 66 169 67
rect 271 67 287 71
rect 267 66 287 67
rect 159 63 169 64
rect 163 59 169 63
rect 267 56 287 64
rect -106 54 -96 55
rect -47 52 -46 56
rect -160 51 -150 52
rect -160 47 -154 51
rect -106 51 -96 52
rect -106 47 -100 51
rect -51 46 -46 52
rect -44 50 -39 56
rect 141 51 157 55
rect 141 50 161 51
rect -44 46 -43 50
rect 267 53 287 54
rect 267 49 283 53
rect 141 40 161 48
rect 141 37 161 38
rect 145 33 161 37
rect -347 5 -342 11
rect -343 1 -342 5
rect -340 7 -338 11
rect -334 7 -332 11
rect -340 1 -332 7
rect -330 5 -325 11
rect -298 6 -292 10
rect -302 5 -292 6
rect -149 6 -143 10
rect -149 5 -139 6
rect -330 1 -329 5
rect -302 1 -292 3
rect -302 -3 -296 1
rect -302 -5 -292 -3
rect -149 1 -139 3
rect 283 26 289 30
rect 279 25 289 26
rect 323 26 324 30
rect 95 15 111 19
rect 279 22 289 23
rect 279 18 285 22
rect 91 14 111 15
rect -145 -3 -139 1
rect -149 -5 -139 -3
rect -66 -2 -65 2
rect -302 -8 -292 -7
rect -343 -14 -342 -10
rect -347 -30 -342 -14
rect -340 -30 -332 -10
rect -330 -26 -325 -10
rect -298 -12 -292 -8
rect -149 -8 -139 -7
rect -70 -8 -65 -2
rect -63 -2 -62 2
rect -63 -8 -58 -2
rect -47 -2 -46 2
rect -51 -8 -46 -2
rect -44 -4 -39 2
rect 91 4 111 12
rect 137 8 143 12
rect 133 7 143 8
rect 286 8 292 12
rect 319 10 324 26
rect 326 10 334 30
rect 336 14 341 30
rect 336 10 337 14
rect 286 7 296 8
rect 133 3 143 5
rect 91 1 111 2
rect 91 -3 107 1
rect 133 -1 139 3
rect 133 -3 143 -1
rect 286 3 296 5
rect 290 -1 296 3
rect 286 -3 296 -1
rect -44 -8 -43 -4
rect -149 -12 -143 -8
rect 9 -9 14 -3
rect 13 -13 14 -9
rect 16 -7 17 -3
rect 323 -5 324 -1
rect 16 -13 21 -7
rect 133 -6 143 -5
rect 137 -10 143 -6
rect 286 -6 296 -5
rect 286 -10 292 -6
rect 319 -11 324 -5
rect 326 -7 334 -1
rect 326 -11 328 -7
rect 332 -11 334 -7
rect 336 -5 337 -1
rect 336 -11 341 -5
rect -291 -22 -285 -18
rect -295 -23 -285 -22
rect -330 -30 -329 -26
rect -295 -26 -285 -25
rect -295 -30 -289 -26
rect 100 -33 105 -27
rect -167 -37 -151 -33
rect 104 -37 105 -33
rect 107 -33 112 -27
rect 107 -37 108 -33
rect 119 -33 124 -27
rect 123 -37 124 -33
rect 126 -31 127 -27
rect 126 -37 131 -31
rect -167 -38 -147 -37
rect -167 -48 -147 -40
rect -289 -53 -273 -49
rect -293 -54 -273 -53
rect -167 -51 -147 -50
rect -163 -55 -147 -51
rect -293 -64 -273 -56
rect 13 -59 14 -55
rect -175 -63 -169 -59
rect -175 -64 -165 -63
rect 9 -65 14 -59
rect 16 -61 24 -55
rect 16 -65 18 -61
rect 22 -65 24 -61
rect 26 -59 27 -55
rect 26 -65 31 -59
rect -293 -67 -273 -66
rect -293 -71 -277 -67
rect -175 -67 -165 -66
rect -171 -71 -165 -67
rect 56 -67 57 -63
rect 52 -83 57 -67
rect 59 -83 67 -63
rect 69 -79 74 -63
rect 69 -83 70 -79
rect -298 -94 -292 -90
rect -302 -95 -292 -94
rect -302 -99 -292 -97
rect -302 -103 -296 -99
rect -302 -105 -292 -103
rect -202 -102 -196 -98
rect -206 -103 -196 -102
rect -148 -102 -142 -98
rect -152 -103 -142 -102
rect -206 -106 -196 -105
rect -302 -108 -292 -107
rect -298 -112 -292 -108
rect -206 -110 -200 -106
rect -152 -106 -142 -105
rect -152 -110 -146 -106
rect -38 -107 -32 -103
rect -42 -108 -32 -107
rect -42 -111 -32 -110
rect -38 -115 -32 -111
rect -291 -122 -285 -118
rect -295 -123 -285 -122
rect -206 -121 -200 -117
rect -206 -122 -196 -121
rect -295 -126 -285 -125
rect -295 -130 -289 -126
rect -206 -125 -196 -124
rect -206 -129 -200 -125
rect -92 -126 -86 -122
rect -96 -127 -86 -126
rect -38 -126 -32 -122
rect 82 -85 83 -81
rect 78 -91 83 -85
rect 85 -87 90 -81
rect 85 -91 86 -87
rect 119 -87 124 -81
rect 123 -91 124 -87
rect 126 -85 127 -81
rect 126 -91 131 -85
rect -42 -127 -32 -126
rect -96 -130 -86 -129
rect -96 -134 -90 -130
rect -42 -130 -32 -129
rect -42 -134 -36 -130
rect 176 -155 181 -149
rect 180 -159 181 -155
rect 183 -153 184 -149
rect 183 -159 188 -153
rect 37 -207 42 -201
rect 9 -214 14 -208
rect 13 -218 14 -214
rect 16 -212 18 -208
rect 22 -212 24 -208
rect 16 -218 24 -212
rect 26 -214 31 -208
rect 41 -211 42 -207
rect 44 -205 45 -201
rect 44 -211 49 -205
rect 68 -205 73 -189
rect 72 -209 73 -205
rect 75 -209 83 -189
rect 85 -193 86 -189
rect 85 -209 90 -193
rect 137 -207 142 -201
rect 26 -218 27 -214
rect 109 -214 114 -208
rect 113 -218 114 -214
rect 116 -212 118 -208
rect 122 -212 124 -208
rect 116 -218 124 -212
rect 126 -214 131 -208
rect 141 -211 142 -207
rect 144 -205 145 -201
rect 144 -211 149 -205
rect 176 -209 181 -203
rect 126 -218 127 -214
rect 180 -213 181 -209
rect 183 -207 184 -203
rect 183 -213 188 -207
rect 199 -207 200 -203
rect 195 -213 200 -207
rect 202 -207 203 -203
rect 202 -213 207 -207
rect 7 -245 13 -241
rect 7 -246 17 -245
rect 28 -245 44 -241
rect 28 -246 48 -245
rect 7 -250 17 -248
rect 11 -254 17 -250
rect 7 -256 17 -254
rect 28 -256 48 -248
rect 7 -259 17 -258
rect 7 -263 13 -259
rect 28 -259 48 -258
rect 32 -263 48 -259
<< pdiffusion >>
rect -48 259 -32 263
rect -52 258 -32 259
rect 48 259 84 263
rect 48 258 88 259
rect -52 254 -32 256
rect -52 250 -36 254
rect -52 248 -32 250
rect 48 248 88 256
rect -52 245 -32 246
rect -48 241 -32 245
rect 48 245 88 246
rect 52 241 88 245
rect -54 214 -53 218
rect -58 198 -53 214
rect -51 202 -43 218
rect -51 198 -49 202
rect -45 198 -43 202
rect -41 214 -40 218
rect -41 198 -36 214
rect -17 183 -12 199
rect -13 179 -12 183
rect -10 195 -9 199
rect -10 179 -5 195
rect 1 183 6 219
rect 5 179 6 183
rect 8 179 16 219
rect 18 215 19 219
rect 18 179 23 215
rect 76 161 81 177
rect 80 157 81 161
rect 83 173 84 177
rect 83 157 88 173
rect 231 152 247 156
rect 227 151 247 152
rect 227 147 247 149
rect -138 139 -122 143
rect -138 138 -118 139
rect -138 135 -118 136
rect -138 131 -122 135
rect 227 143 243 147
rect 227 141 247 143
rect 227 138 247 139
rect 231 134 247 138
rect -193 120 -177 124
rect -193 119 -173 120
rect -138 120 -122 124
rect -138 119 -118 120
rect 165 130 181 134
rect 161 129 181 130
rect 161 126 181 127
rect 161 122 177 126
rect -193 116 -173 117
rect -189 112 -173 116
rect -138 116 -118 117
rect -134 112 -118 116
rect 57 106 62 122
rect 61 102 62 106
rect 64 106 69 122
rect 64 102 65 106
rect 76 106 81 122
rect 80 102 81 106
rect 83 118 84 122
rect 83 102 88 118
rect 165 112 201 116
rect 161 111 201 112
rect 161 101 201 109
rect 227 108 263 112
rect 227 107 267 108
rect 161 98 201 99
rect 161 94 197 98
rect 227 97 267 105
rect 227 94 267 95
rect 231 90 267 94
rect -138 74 -122 78
rect -138 73 -118 74
rect -51 73 -46 89
rect -347 34 -342 70
rect -343 30 -342 34
rect -340 30 -332 70
rect -330 34 -325 70
rect -138 70 -118 71
rect -138 66 -122 70
rect -47 69 -46 73
rect -44 85 -43 89
rect -44 69 -39 85
rect -193 55 -177 59
rect -193 54 -173 55
rect -138 55 -122 59
rect -138 54 -118 55
rect 185 67 201 71
rect 181 66 201 67
rect 231 67 247 71
rect 227 66 247 67
rect 323 66 324 70
rect 181 63 201 64
rect 181 59 197 63
rect 227 62 247 64
rect 227 58 243 62
rect 227 56 247 58
rect -193 51 -173 52
rect -189 47 -173 51
rect -138 51 -118 52
rect -134 47 -118 51
rect 181 51 197 55
rect 181 50 201 51
rect 227 53 247 54
rect 231 49 247 53
rect 319 50 324 66
rect 326 54 334 70
rect 326 50 328 54
rect 332 50 334 54
rect 336 66 337 70
rect 336 50 341 66
rect 181 46 201 48
rect 185 42 201 46
rect 181 40 201 42
rect -330 30 -329 34
rect -70 18 -65 34
rect -66 14 -65 18
rect -63 18 -58 34
rect -63 14 -62 18
rect -51 18 -46 34
rect -47 14 -46 18
rect -44 30 -43 34
rect 181 37 201 38
rect 181 33 197 37
rect -44 14 -39 30
rect 13 25 14 29
rect -273 6 -237 10
rect -273 5 -233 6
rect -204 6 -168 10
rect -208 5 -168 6
rect -273 -5 -233 3
rect -208 -5 -168 3
rect 9 9 14 25
rect 16 13 21 29
rect 247 26 263 30
rect 247 25 267 26
rect 247 22 267 23
rect 55 15 71 19
rect 51 14 71 15
rect 251 18 267 22
rect 16 9 17 13
rect 51 10 71 12
rect -273 -8 -233 -7
rect -269 -12 -233 -8
rect -208 -8 -168 -7
rect -208 -12 -172 -8
rect 51 6 67 10
rect 51 4 71 6
rect 166 8 202 12
rect 162 7 202 8
rect 227 8 263 12
rect 227 7 267 8
rect 51 1 71 2
rect 55 -3 71 1
rect 162 -3 202 5
rect 227 -3 267 5
rect 162 -6 202 -5
rect 162 -10 176 -6
rect 180 -10 198 -6
rect 227 -6 267 -5
rect 231 -10 267 -6
rect -273 -22 -257 -18
rect -273 -23 -253 -22
rect -273 -26 -253 -25
rect -269 -30 -253 -26
rect -203 -37 -187 -33
rect -207 -38 -187 -37
rect 323 -34 324 -30
rect -207 -42 -187 -40
rect -207 -46 -191 -42
rect -207 -48 -187 -46
rect -347 -66 -342 -50
rect -343 -70 -342 -66
rect -340 -54 -338 -50
rect -334 -54 -332 -50
rect -340 -70 -332 -54
rect -330 -66 -325 -50
rect -253 -53 -237 -49
rect -253 -54 -233 -53
rect -207 -51 -187 -50
rect -203 -55 -187 -51
rect 104 -53 105 -49
rect -253 -58 -233 -56
rect -249 -62 -233 -58
rect -253 -64 -233 -62
rect -203 -63 -187 -59
rect -207 -64 -187 -63
rect -330 -70 -329 -66
rect -253 -67 -233 -66
rect -253 -71 -237 -67
rect -207 -67 -187 -66
rect -207 -71 -191 -67
rect 100 -69 105 -53
rect 107 -53 108 -49
rect 107 -69 112 -53
rect 123 -53 124 -49
rect 119 -69 124 -53
rect 126 -65 131 -49
rect 126 -69 127 -65
rect 319 -70 324 -34
rect 326 -70 334 -30
rect 336 -34 337 -30
rect 336 -70 341 -34
rect -273 -94 -237 -90
rect -273 -95 -233 -94
rect -273 -105 -233 -97
rect -184 -102 -168 -98
rect -184 -103 -164 -102
rect -129 -102 -113 -98
rect -129 -103 -109 -102
rect -273 -108 -233 -107
rect -269 -112 -233 -108
rect -184 -106 -164 -105
rect -180 -110 -164 -106
rect -129 -106 -109 -105
rect -125 -110 -109 -106
rect -74 -107 -58 -103
rect -74 -108 -54 -107
rect -74 -111 -54 -110
rect -74 -115 -58 -111
rect -273 -122 -257 -118
rect -180 -121 -164 -117
rect -184 -122 -164 -121
rect 9 -120 14 -84
rect -273 -123 -253 -122
rect -273 -126 -253 -125
rect -269 -130 -253 -126
rect -184 -125 -164 -124
rect -180 -129 -164 -125
rect -129 -126 -113 -122
rect -129 -127 -109 -126
rect -74 -126 -58 -122
rect -74 -127 -54 -126
rect 13 -124 14 -120
rect 16 -124 24 -84
rect 26 -88 27 -84
rect 26 -124 31 -88
rect 52 -119 57 -103
rect 56 -123 57 -119
rect 59 -107 61 -103
rect 65 -107 67 -103
rect 59 -123 67 -107
rect 69 -119 74 -103
rect 69 -123 70 -119
rect 78 -119 83 -103
rect 82 -123 83 -119
rect 85 -107 86 -103
rect 85 -123 90 -107
rect 123 -108 124 -104
rect 119 -124 124 -108
rect 126 -120 131 -104
rect 126 -124 127 -120
rect 180 -120 181 -116
rect -129 -130 -109 -129
rect -125 -134 -109 -130
rect -74 -130 -54 -129
rect -70 -134 -54 -130
rect 176 -136 181 -120
rect 183 -132 188 -116
rect 183 -136 184 -132
rect 13 -153 14 -149
rect 9 -189 14 -153
rect 16 -189 24 -149
rect 26 -185 31 -149
rect 72 -153 73 -149
rect 68 -169 73 -153
rect 75 -165 83 -149
rect 75 -169 77 -165
rect 81 -169 83 -165
rect 85 -153 86 -149
rect 85 -169 90 -153
rect 113 -153 114 -149
rect 26 -189 27 -185
rect 41 -173 42 -169
rect 37 -189 42 -173
rect 44 -185 49 -169
rect 44 -189 45 -185
rect 109 -189 114 -153
rect 116 -189 124 -149
rect 126 -185 131 -149
rect 126 -189 127 -185
rect 141 -173 142 -169
rect 137 -189 142 -173
rect 144 -185 149 -169
rect 144 -189 145 -185
rect 180 -175 181 -171
rect 176 -191 181 -175
rect 183 -187 188 -171
rect 183 -191 184 -187
rect 195 -187 200 -171
rect 199 -191 200 -187
rect 202 -187 207 -171
rect 202 -191 203 -187
rect -52 -245 -16 -241
rect -52 -246 -12 -245
rect 68 -245 84 -241
rect 68 -246 88 -245
rect -52 -256 -12 -248
rect 68 -250 88 -248
rect 72 -254 88 -250
rect 68 -256 88 -254
rect -52 -259 -12 -258
rect -52 -263 -16 -259
rect 68 -259 88 -258
rect 68 -263 84 -259
<< ndcontact >>
rect 4 259 8 263
rect 19 259 23 263
rect 25 250 29 254
rect -12 241 -8 245
rect 19 241 23 245
rect -58 174 -54 178
rect -40 158 -36 162
rect -17 163 -13 167
rect -9 157 -5 161
rect 1 150 5 154
rect 10 156 14 160
rect 19 150 23 154
rect 267 152 271 156
rect -106 139 -102 143
rect 76 140 80 144
rect -106 131 -102 135
rect 84 134 88 138
rect 283 134 287 138
rect -160 120 -156 124
rect -106 120 -102 124
rect 145 130 149 134
rect 139 122 143 126
rect -154 112 -150 116
rect -100 112 -96 116
rect 132 112 136 116
rect 138 103 142 107
rect 292 108 296 112
rect 132 94 136 98
rect 286 99 290 103
rect 292 90 296 94
rect -106 74 -102 78
rect -106 66 -102 70
rect 57 86 61 90
rect 65 86 69 90
rect 76 86 80 90
rect 84 80 88 84
rect -160 55 -156 59
rect -106 55 -102 59
rect 165 67 169 71
rect 267 67 271 71
rect 159 59 163 63
rect -51 52 -47 56
rect -154 47 -150 51
rect -100 47 -96 51
rect 157 51 161 55
rect -43 46 -39 50
rect 283 49 287 53
rect 141 33 145 37
rect -347 1 -343 5
rect -338 7 -334 11
rect -302 6 -298 10
rect -143 6 -139 10
rect -329 1 -325 5
rect -296 -3 -292 1
rect 279 26 283 30
rect 319 26 323 30
rect 91 15 95 19
rect 285 18 289 22
rect -149 -3 -145 1
rect -70 -2 -66 2
rect -347 -14 -343 -10
rect -302 -12 -298 -8
rect -62 -2 -58 2
rect -51 -2 -47 2
rect 133 8 137 12
rect 292 8 296 12
rect 337 10 341 14
rect 107 -3 111 1
rect 139 -1 143 3
rect 286 -1 290 3
rect -43 -8 -39 -4
rect -143 -12 -139 -8
rect 9 -13 13 -9
rect 17 -7 21 -3
rect 319 -5 323 -1
rect 133 -10 137 -6
rect 292 -10 296 -6
rect 328 -11 332 -7
rect 337 -5 341 -1
rect -295 -22 -291 -18
rect -329 -30 -325 -26
rect -289 -30 -285 -26
rect -151 -37 -147 -33
rect 100 -37 104 -33
rect 108 -37 112 -33
rect 119 -37 123 -33
rect 127 -31 131 -27
rect -293 -53 -289 -49
rect -167 -55 -163 -51
rect 9 -59 13 -55
rect -169 -63 -165 -59
rect 18 -65 22 -61
rect 27 -59 31 -55
rect -277 -71 -273 -67
rect -175 -71 -171 -67
rect 52 -67 56 -63
rect 70 -83 74 -79
rect -302 -94 -298 -90
rect -296 -103 -292 -99
rect -206 -102 -202 -98
rect -152 -102 -148 -98
rect -302 -112 -298 -108
rect -200 -110 -196 -106
rect -146 -110 -142 -106
rect -42 -107 -38 -103
rect -42 -115 -38 -111
rect -295 -122 -291 -118
rect -200 -121 -196 -117
rect -289 -130 -285 -126
rect -200 -129 -196 -125
rect -96 -126 -92 -122
rect -42 -126 -38 -122
rect 78 -85 82 -81
rect 86 -91 90 -87
rect 119 -91 123 -87
rect 127 -85 131 -81
rect -90 -134 -86 -130
rect -36 -134 -32 -130
rect 176 -159 180 -155
rect 184 -153 188 -149
rect 9 -218 13 -214
rect 18 -212 22 -208
rect 37 -211 41 -207
rect 45 -205 49 -201
rect 68 -209 72 -205
rect 86 -193 90 -189
rect 27 -218 31 -214
rect 109 -218 113 -214
rect 118 -212 122 -208
rect 137 -211 141 -207
rect 145 -205 149 -201
rect 127 -218 131 -214
rect 176 -213 180 -209
rect 184 -207 188 -203
rect 195 -207 199 -203
rect 203 -207 207 -203
rect 13 -245 17 -241
rect 44 -245 48 -241
rect 7 -254 11 -250
rect 13 -263 17 -259
rect 28 -263 32 -259
<< pdcontact >>
rect -52 259 -48 263
rect 84 259 88 263
rect -36 250 -32 254
rect -52 241 -48 245
rect 48 241 52 245
rect -58 214 -54 218
rect -49 198 -45 202
rect -40 214 -36 218
rect -17 179 -13 183
rect -9 195 -5 199
rect 1 179 5 183
rect 19 215 23 219
rect 76 157 80 161
rect 84 173 88 177
rect 227 152 231 156
rect -122 139 -118 143
rect -122 131 -118 135
rect 243 143 247 147
rect 227 134 231 138
rect -177 120 -173 124
rect -122 120 -118 124
rect 161 130 165 134
rect 177 122 181 126
rect -193 112 -189 116
rect -138 112 -134 116
rect 57 102 61 106
rect 65 102 69 106
rect 76 102 80 106
rect 84 118 88 122
rect 161 112 165 116
rect 263 108 267 112
rect 197 94 201 98
rect 227 90 231 94
rect -122 74 -118 78
rect -347 30 -343 34
rect -122 66 -118 70
rect -51 69 -47 73
rect -43 85 -39 89
rect -177 55 -173 59
rect -122 55 -118 59
rect 181 67 185 71
rect 227 67 231 71
rect 319 66 323 70
rect 197 59 201 63
rect 243 58 247 62
rect -193 47 -189 51
rect -138 47 -134 51
rect 197 51 201 55
rect 227 49 231 53
rect 328 50 332 54
rect 337 66 341 70
rect 181 42 185 46
rect -329 30 -325 34
rect -70 14 -66 18
rect -62 14 -58 18
rect -51 14 -47 18
rect -43 30 -39 34
rect 197 33 201 37
rect 9 25 13 29
rect -237 6 -233 10
rect -208 6 -204 10
rect 263 26 267 30
rect 51 15 55 19
rect 247 18 251 22
rect 17 9 21 13
rect -273 -12 -269 -8
rect -172 -12 -168 -8
rect 67 6 71 10
rect 162 8 166 12
rect 263 8 267 12
rect 51 -3 55 1
rect 176 -10 180 -6
rect 198 -10 202 -6
rect 227 -10 231 -6
rect -257 -22 -253 -18
rect -273 -30 -269 -26
rect -207 -37 -203 -33
rect 319 -34 323 -30
rect -191 -46 -187 -42
rect -347 -70 -343 -66
rect -338 -54 -334 -50
rect -237 -53 -233 -49
rect -207 -55 -203 -51
rect 100 -53 104 -49
rect -253 -62 -249 -58
rect -207 -63 -203 -59
rect -329 -70 -325 -66
rect -237 -71 -233 -67
rect -191 -71 -187 -67
rect 108 -53 112 -49
rect 119 -53 123 -49
rect 127 -69 131 -65
rect 337 -34 341 -30
rect -237 -94 -233 -90
rect -168 -102 -164 -98
rect -113 -102 -109 -98
rect -273 -112 -269 -108
rect -184 -110 -180 -106
rect -129 -110 -125 -106
rect -58 -107 -54 -103
rect -58 -115 -54 -111
rect -257 -122 -253 -118
rect -184 -121 -180 -117
rect -273 -130 -269 -126
rect -184 -129 -180 -125
rect -113 -126 -109 -122
rect -58 -126 -54 -122
rect 9 -124 13 -120
rect 27 -88 31 -84
rect 52 -123 56 -119
rect 61 -107 65 -103
rect 70 -123 74 -119
rect 78 -123 82 -119
rect 86 -107 90 -103
rect 119 -108 123 -104
rect 127 -124 131 -120
rect 176 -120 180 -116
rect -129 -134 -125 -130
rect -74 -134 -70 -130
rect 184 -136 188 -132
rect 9 -153 13 -149
rect 68 -153 72 -149
rect 77 -169 81 -165
rect 86 -153 90 -149
rect 109 -153 113 -149
rect 27 -189 31 -185
rect 37 -173 41 -169
rect 45 -189 49 -185
rect 127 -189 131 -185
rect 137 -173 141 -169
rect 145 -189 149 -185
rect 176 -175 180 -171
rect 184 -191 188 -187
rect 195 -191 199 -187
rect 203 -191 207 -187
rect -16 -245 -12 -241
rect 84 -245 88 -241
rect 68 -254 72 -250
rect -16 -263 -12 -259
rect 84 -263 88 -259
<< polysilicon >>
rect -56 256 -52 258
rect -32 256 -12 258
rect 8 256 11 258
rect 16 256 19 258
rect 29 256 48 258
rect 88 256 91 258
rect -56 246 -52 248
rect -32 246 -12 248
rect 8 246 11 248
rect 16 246 19 248
rect 29 246 48 248
rect 88 246 91 248
rect -53 218 -51 222
rect -43 218 -41 222
rect 6 219 8 222
rect 16 219 18 222
rect -12 199 -10 203
rect -53 178 -51 198
rect -43 178 -41 198
rect -12 167 -10 179
rect -53 155 -51 158
rect -43 155 -41 158
rect 6 160 8 179
rect 16 160 18 179
rect 81 177 83 181
rect -12 153 -10 157
rect 6 147 8 150
rect 16 147 18 150
rect 81 144 83 157
rect 223 149 227 151
rect 247 149 267 151
rect 287 149 290 151
rect -150 136 -138 138
rect -118 136 -115 138
rect -109 136 -106 138
rect -96 136 -90 138
rect 223 139 227 141
rect 247 139 267 141
rect 287 139 290 141
rect 62 122 64 134
rect 81 130 83 134
rect 135 127 139 129
rect 149 127 161 129
rect 181 127 185 129
rect 81 122 83 126
rect -197 117 -193 119
rect -173 117 -160 119
rect -150 117 -146 119
rect -142 117 -138 119
rect -118 117 -106 119
rect -96 117 -93 119
rect 129 109 132 111
rect 142 109 161 111
rect 201 109 204 111
rect 62 99 64 102
rect -46 89 -44 93
rect 62 90 64 93
rect 81 90 83 102
rect 224 105 227 107
rect 267 105 286 107
rect 296 105 299 107
rect 129 99 132 101
rect 142 99 161 101
rect 201 99 204 101
rect 224 95 227 97
rect 267 95 286 97
rect 296 95 299 97
rect -342 70 -340 73
rect -332 70 -330 73
rect -150 71 -138 73
rect -118 71 -115 73
rect -109 71 -106 73
rect -96 71 -90 73
rect 62 74 64 80
rect 81 77 83 80
rect -46 56 -44 69
rect 324 70 326 74
rect 334 70 336 74
rect 155 64 159 66
rect 169 64 181 66
rect 201 64 205 66
rect 223 64 227 66
rect 247 64 267 66
rect 287 64 290 66
rect -197 52 -193 54
rect -173 52 -160 54
rect -150 52 -146 54
rect -142 52 -138 54
rect -118 52 -106 54
rect -96 52 -93 54
rect 223 54 227 56
rect 247 54 267 56
rect 287 54 290 56
rect 138 48 141 50
rect 161 48 181 50
rect 201 48 205 50
rect -65 34 -63 46
rect -46 42 -44 46
rect 138 38 141 40
rect 161 38 181 40
rect 201 38 205 40
rect -46 34 -44 38
rect -342 11 -340 30
rect -332 11 -330 30
rect 14 29 16 33
rect 324 30 326 50
rect 334 30 336 50
rect -65 11 -63 14
rect -305 3 -302 5
rect -292 3 -273 5
rect -233 3 -230 5
rect -211 3 -208 5
rect -168 3 -149 5
rect -139 3 -136 5
rect -342 -2 -340 1
rect -332 -2 -330 1
rect -65 2 -63 5
rect -46 2 -44 14
rect 243 23 247 25
rect 267 23 279 25
rect 289 23 293 25
rect 47 12 51 14
rect 71 12 91 14
rect 111 12 114 14
rect -305 -7 -302 -5
rect -292 -7 -273 -5
rect -233 -7 -230 -5
rect -211 -7 -208 -5
rect -168 -7 -149 -5
rect -139 -7 -136 -5
rect -342 -10 -340 -7
rect -332 -10 -330 -7
rect 14 -3 16 9
rect 324 7 326 10
rect 334 7 336 10
rect 130 5 133 7
rect 143 5 162 7
rect 202 5 205 7
rect 224 5 227 7
rect 267 5 286 7
rect 296 5 299 7
rect 47 2 51 4
rect 71 2 91 4
rect 111 2 114 4
rect 324 -1 326 2
rect 334 -1 336 2
rect -65 -14 -63 -8
rect -46 -11 -44 -8
rect 130 -5 133 -3
rect 143 -5 162 -3
rect 202 -5 205 -3
rect 224 -5 227 -3
rect 267 -5 286 -3
rect 296 -5 299 -3
rect 14 -17 16 -13
rect -299 -25 -295 -23
rect -285 -25 -273 -23
rect -253 -25 -249 -23
rect 105 -27 107 -21
rect 124 -27 126 -24
rect -342 -50 -340 -30
rect -332 -50 -330 -30
rect 324 -30 326 -11
rect 334 -30 336 -11
rect -211 -40 -207 -38
rect -187 -40 -167 -38
rect -147 -40 -144 -38
rect 105 -40 107 -37
rect -211 -50 -207 -48
rect -187 -50 -167 -48
rect -147 -50 -144 -48
rect 105 -49 107 -46
rect 124 -49 126 -37
rect -296 -56 -293 -54
rect -273 -56 -253 -54
rect -233 -56 -229 -54
rect 14 -55 16 -52
rect 24 -55 26 -52
rect -296 -66 -293 -64
rect -273 -66 -253 -64
rect -233 -66 -229 -64
rect -211 -66 -207 -64
rect -187 -66 -175 -64
rect -165 -66 -161 -64
rect 57 -63 59 -60
rect 67 -63 69 -60
rect -342 -74 -340 -70
rect -332 -74 -330 -70
rect 14 -84 16 -65
rect 24 -84 26 -65
rect 83 -81 85 -77
rect 105 -81 107 -69
rect 124 -73 126 -69
rect 324 -73 326 -70
rect 334 -73 336 -70
rect 124 -81 126 -77
rect -305 -97 -302 -95
rect -292 -97 -273 -95
rect -233 -97 -230 -95
rect -209 -105 -206 -103
rect -196 -105 -184 -103
rect -164 -105 -160 -103
rect -156 -105 -152 -103
rect -142 -105 -129 -103
rect -109 -105 -105 -103
rect -305 -107 -302 -105
rect -292 -107 -273 -105
rect -233 -107 -230 -105
rect -86 -110 -74 -108
rect -54 -110 -51 -108
rect -45 -110 -42 -108
rect -32 -110 -26 -108
rect -299 -125 -295 -123
rect -285 -125 -273 -123
rect -253 -125 -249 -123
rect -212 -124 -206 -122
rect -196 -124 -193 -122
rect -187 -124 -184 -122
rect -164 -124 -152 -122
rect 57 -103 59 -83
rect 67 -103 69 -83
rect 83 -103 85 -91
rect 124 -104 126 -91
rect 14 -127 16 -124
rect 24 -127 26 -124
rect 57 -127 59 -123
rect 67 -127 69 -123
rect 83 -127 85 -123
rect 181 -116 183 -112
rect -133 -129 -129 -127
rect -109 -129 -96 -127
rect -86 -129 -82 -127
rect -78 -129 -74 -127
rect -54 -129 -42 -127
rect -32 -129 -29 -127
rect 124 -128 126 -124
rect 14 -149 16 -146
rect 24 -149 26 -146
rect 73 -149 75 -145
rect 83 -149 85 -145
rect 114 -149 116 -146
rect 124 -149 126 -146
rect 181 -149 183 -136
rect 42 -169 44 -165
rect 73 -189 75 -169
rect 83 -189 85 -169
rect 181 -163 183 -159
rect 142 -169 144 -165
rect 181 -171 183 -167
rect 200 -171 202 -159
rect 14 -208 16 -189
rect 24 -208 26 -189
rect 42 -201 44 -189
rect 114 -208 116 -189
rect 124 -208 126 -189
rect 142 -201 144 -189
rect 42 -215 44 -211
rect 73 -212 75 -209
rect 83 -212 85 -209
rect 181 -203 183 -191
rect 200 -194 202 -191
rect 200 -203 202 -200
rect 142 -215 144 -211
rect 181 -216 183 -213
rect 14 -221 16 -218
rect 24 -221 26 -218
rect 114 -221 116 -218
rect 124 -221 126 -218
rect 200 -219 202 -213
rect -55 -248 -52 -246
rect -12 -248 7 -246
rect 17 -248 20 -246
rect 25 -248 28 -246
rect 48 -248 68 -246
rect 88 -248 92 -246
rect -55 -258 -52 -256
rect -12 -258 7 -256
rect 17 -258 20 -256
rect 25 -258 28 -256
rect 48 -258 68 -256
rect 88 -258 92 -256
<< polycontact >>
rect -25 258 -21 262
rect 30 258 34 262
rect -17 248 -13 252
rect 37 248 41 252
rect -51 179 -47 183
rect -41 187 -37 191
rect -10 168 -6 172
rect 8 168 12 172
rect 18 161 22 165
rect 83 145 87 149
rect -95 138 -91 142
rect -149 132 -145 136
rect 262 145 266 149
rect 254 135 258 139
rect 64 129 68 133
rect 150 123 154 127
rect -165 113 -161 117
rect -111 113 -107 117
rect 150 105 154 109
rect 83 91 87 95
rect 143 95 147 99
rect 274 101 278 105
rect 281 91 285 95
rect -95 73 -91 77
rect -149 67 -145 71
rect 58 75 62 79
rect -44 57 -40 61
rect 170 60 174 64
rect 262 60 266 64
rect -165 48 -161 52
rect -111 48 -107 52
rect 254 50 258 54
rect -63 41 -59 45
rect 162 44 166 48
rect -346 12 -342 16
rect -336 19 -332 23
rect 170 34 174 38
rect 326 31 330 35
rect 336 39 340 43
rect -291 5 -287 9
rect -154 5 -150 9
rect -284 -5 -280 -1
rect 274 19 278 23
rect -44 3 -40 7
rect -161 -5 -157 -1
rect 10 -2 14 2
rect 86 8 90 12
rect 78 -2 82 2
rect 151 1 155 5
rect 274 1 278 5
rect -69 -13 -65 -9
rect 144 -9 148 -5
rect 281 -9 285 -5
rect -284 -23 -280 -19
rect 101 -26 105 -22
rect -346 -43 -342 -39
rect -336 -35 -332 -31
rect -180 -38 -176 -34
rect 326 -23 330 -19
rect 336 -16 340 -12
rect -172 -48 -168 -44
rect -264 -54 -260 -50
rect 126 -42 130 -38
rect -272 -64 -268 -60
rect -180 -64 -176 -60
rect 10 -70 14 -66
rect 20 -77 24 -73
rect 107 -80 111 -76
rect -291 -95 -287 -91
rect -284 -105 -280 -101
rect -195 -103 -191 -99
rect -141 -103 -137 -99
rect -31 -108 -27 -104
rect -85 -114 -81 -110
rect -284 -123 -280 -119
rect -157 -122 -153 -118
rect -211 -128 -207 -124
rect 53 -96 57 -92
rect 63 -88 67 -84
rect 79 -96 83 -92
rect 126 -96 130 -92
rect -101 -133 -97 -129
rect -47 -133 -43 -129
rect 177 -148 181 -144
rect 69 -180 73 -176
rect 79 -188 83 -184
rect 196 -164 200 -160
rect 10 -207 14 -203
rect 20 -200 24 -196
rect 38 -200 42 -196
rect 110 -207 114 -203
rect 120 -200 124 -196
rect 138 -200 142 -196
rect 177 -202 181 -198
rect 202 -218 206 -214
rect -5 -252 -1 -248
rect 49 -252 53 -248
rect 2 -262 6 -258
rect 57 -262 61 -258
<< metal1 >>
rect -62 290 98 293
rect -62 263 -59 290
rect -6 283 -3 287
rect -25 275 41 278
rect -62 259 -52 263
rect -25 262 -21 275
rect -62 246 -59 259
rect -17 269 20 272
rect -32 250 -21 254
rect -25 245 -21 250
rect -17 252 -13 269
rect 25 269 34 272
rect 8 259 19 263
rect 30 262 34 269
rect 12 245 15 259
rect 29 250 34 254
rect 30 245 34 250
rect 37 252 41 275
rect 95 263 98 290
rect 88 259 116 263
rect -59 241 -52 245
rect -25 241 -12 245
rect 12 244 19 245
rect -25 234 -21 241
rect 16 241 19 244
rect 30 241 48 245
rect 30 235 34 241
rect -93 231 -21 234
rect -93 164 -90 231
rect -70 227 -36 228
rect -67 225 -36 227
rect -58 218 -54 225
rect -40 218 -36 225
rect -49 191 -45 198
rect -28 191 -25 231
rect 94 231 111 234
rect -9 226 23 229
rect -9 199 -5 226
rect 19 219 23 226
rect 37 225 87 228
rect 37 219 40 225
rect 23 215 40 219
rect -172 161 -90 164
rect -87 188 -45 191
rect -172 134 -169 161
rect -87 155 -84 188
rect -111 152 -84 155
rect -111 143 -107 152
rect -118 139 -106 143
rect -95 142 -91 144
rect -209 131 -169 134
rect -209 35 -206 131
rect -149 130 -145 132
rect -118 131 -106 135
rect -111 130 -106 131
rect -95 130 -91 138
rect -111 124 -106 125
rect -173 120 -160 124
rect -118 120 -106 124
rect -375 30 -347 34
rect -375 -77 -372 30
rect -362 19 -336 23
rect -362 -39 -359 19
rect -329 16 -325 30
rect -284 32 -206 35
rect -203 112 -193 116
rect -203 51 -200 112
rect -165 105 -161 113
rect -154 97 -150 112
rect -138 105 -134 112
rect -111 108 -107 113
rect -96 112 -95 116
rect -87 108 -84 152
rect -64 150 -61 188
rect -58 178 -54 188
rect -37 187 -25 191
rect 84 189 87 225
rect 108 203 111 231
rect 108 198 168 203
rect -47 179 -27 183
rect -30 172 -27 179
rect -17 172 -13 179
rect 1 172 5 179
rect 84 177 88 184
rect -30 168 -13 172
rect -6 168 5 172
rect 12 168 30 172
rect -17 167 -13 168
rect 1 165 5 168
rect 1 161 14 165
rect 22 161 31 165
rect -40 156 -36 158
rect -40 153 -23 156
rect -9 156 -5 157
rect 10 160 14 161
rect -18 153 -5 156
rect -64 147 -12 150
rect -15 140 -12 147
rect -9 146 -5 153
rect 1 146 5 150
rect 19 146 23 150
rect -9 143 23 146
rect -111 105 -84 108
rect -154 94 -78 97
rect -111 87 -84 90
rect -111 78 -107 87
rect -118 74 -106 78
rect -95 77 -91 79
rect -149 65 -145 67
rect -118 66 -106 70
rect -111 65 -106 66
rect -95 65 -91 73
rect -111 59 -106 60
rect -173 55 -160 59
rect -118 55 -106 59
rect -203 47 -193 51
rect -356 12 -346 16
rect -338 12 -317 16
rect -312 13 -287 16
rect -356 7 -353 12
rect -338 11 -334 12
rect -309 6 -302 10
rect -291 9 -287 13
rect -356 -31 -353 2
rect -347 -3 -343 1
rect -329 -3 -325 1
rect -309 -3 -306 6
rect -292 -3 -287 1
rect -347 -6 -306 -3
rect -347 -10 -343 -6
rect -309 -8 -306 -6
rect -291 -8 -287 -3
rect -284 -1 -281 32
rect -203 24 -200 47
rect -165 40 -161 48
rect -154 29 -150 47
rect -138 40 -134 47
rect -111 44 -107 48
rect -96 47 -95 51
rect -87 43 -84 87
rect -106 40 -84 43
rect -81 29 -78 94
rect -43 89 -39 96
rect -51 56 -47 69
rect -40 57 -32 61
rect -7 57 -4 143
rect -23 54 -4 57
rect 28 64 31 161
rect 76 144 80 157
rect 87 145 95 149
rect 108 138 111 198
rect 123 184 168 189
rect 254 156 258 162
rect 217 152 227 156
rect 254 152 267 156
rect 217 150 220 152
rect 254 147 258 152
rect 150 141 211 144
rect 88 134 128 138
rect 150 134 154 141
rect 68 129 70 133
rect 125 126 128 134
rect 149 130 161 134
rect 208 132 211 141
rect 217 138 220 145
rect 247 143 258 147
rect 217 135 227 138
rect 208 129 217 132
rect 214 127 217 129
rect 254 127 258 135
rect 125 122 139 126
rect 88 118 95 122
rect 125 116 128 122
rect 150 116 154 123
rect 181 122 211 126
rect 214 124 258 127
rect 125 112 132 116
rect 143 112 161 116
rect 57 95 61 102
rect 45 91 61 95
rect 45 71 48 91
rect 57 90 61 91
rect 65 95 69 102
rect 76 95 80 102
rect 125 98 128 112
rect 143 107 147 112
rect 142 103 147 107
rect 65 90 70 95
rect 75 90 80 95
rect 87 91 92 95
rect 128 94 132 98
rect 84 79 88 80
rect 56 75 58 79
rect 62 75 70 79
rect 92 71 95 90
rect 45 68 95 71
rect 143 69 147 95
rect 150 87 154 105
rect 208 98 211 122
rect 262 123 266 145
rect 287 134 300 138
rect 262 120 278 123
rect 274 112 278 120
rect 297 112 300 134
rect 267 108 285 112
rect 296 108 303 112
rect 201 94 208 98
rect 213 94 220 96
rect 213 93 227 94
rect 217 90 227 93
rect 274 83 278 101
rect 281 103 285 108
rect 281 99 286 103
rect 170 80 278 83
rect 300 94 303 108
rect 170 71 174 80
rect 281 77 285 91
rect 296 90 303 94
rect 259 74 285 77
rect 254 71 259 72
rect 128 66 147 69
rect 169 67 181 71
rect 217 67 227 71
rect 254 67 267 71
rect 128 64 131 66
rect 28 61 131 64
rect -23 52 -20 54
rect -39 47 -25 50
rect -39 46 -20 47
rect -59 41 -57 45
rect -39 30 -32 34
rect 9 29 13 49
rect -154 26 -78 29
rect -226 21 -200 24
rect -226 10 -223 21
rect -233 6 -208 10
rect -309 -12 -302 -8
rect -291 -12 -273 -8
rect -309 -18 -306 -12
rect -309 -22 -302 -18
rect -297 -22 -295 -18
rect -284 -19 -280 -12
rect -226 -18 -223 6
rect -253 -22 -223 -18
rect -285 -30 -273 -26
rect -356 -35 -336 -31
rect -329 -39 -325 -30
rect -284 -37 -280 -30
rect -217 -33 -214 6
rect -161 -1 -157 16
rect -153 13 -152 16
rect -154 9 -150 13
rect -138 10 -135 26
rect -139 6 -132 10
rect -70 7 -66 14
rect -154 -3 -149 1
rect -154 -8 -150 -3
rect -135 -8 -132 6
rect -82 3 -66 7
rect -168 -12 -150 -8
rect -139 -12 -136 -8
rect -154 -17 -150 -12
rect -180 -22 -155 -19
rect -82 -17 -79 3
rect -70 2 -66 3
rect -62 7 -58 14
rect -51 7 -47 14
rect -62 2 -57 7
rect -52 2 -47 7
rect -40 3 -32 7
rect -35 2 -32 3
rect 17 2 21 9
rect 28 2 31 61
rect 134 59 159 63
rect 44 39 47 53
rect -35 -1 10 2
rect -43 -9 -39 -8
rect -71 -13 -69 -9
rect -65 -13 -57 -9
rect -35 -17 -32 -1
rect -82 -20 -32 -17
rect -2 -2 10 -1
rect 17 -2 31 2
rect 34 36 47 39
rect -217 -37 -207 -33
rect -180 -34 -176 -22
rect -2 -25 1 -2
rect 17 -3 21 -2
rect -362 -43 -346 -39
rect -338 -43 -318 -39
rect -338 -50 -334 -43
rect -284 -40 -260 -37
rect -313 -43 -287 -40
rect -290 -46 -268 -43
rect -306 -53 -302 -49
rect -297 -53 -293 -49
rect -347 -77 -343 -70
rect -329 -77 -325 -70
rect -375 -80 -330 -77
rect -306 -90 -303 -53
rect -272 -60 -268 -46
rect -264 -50 -260 -40
rect -233 -53 -223 -49
rect -226 -56 -223 -53
rect -217 -51 -214 -37
rect -172 -28 1 -25
rect -187 -46 -176 -42
rect -180 -51 -176 -46
rect -172 -44 -168 -28
rect -147 -37 -143 -33
rect -217 -55 -207 -51
rect -180 -55 -167 -51
rect -217 -56 -214 -55
rect -264 -62 -253 -58
rect -214 -61 -207 -59
rect -264 -67 -260 -62
rect -226 -67 -223 -61
rect -217 -63 -207 -61
rect -180 -60 -176 -55
rect -143 -59 -140 -37
rect -123 -37 -5 -34
rect 9 -48 13 -13
rect 34 -40 37 36
rect 41 19 44 26
rect 78 19 82 50
rect 134 38 137 59
rect 170 55 174 60
rect 201 59 208 63
rect 208 55 211 59
rect 161 51 174 55
rect 201 52 211 55
rect 217 53 220 67
rect 254 62 258 67
rect 247 58 258 62
rect 217 52 227 53
rect 201 51 227 52
rect 138 33 141 37
rect 162 28 166 44
rect 170 46 174 51
rect 208 49 227 51
rect 170 42 181 46
rect 131 25 166 28
rect 208 37 211 44
rect 170 22 174 34
rect 201 33 211 37
rect 144 19 174 22
rect 217 22 220 49
rect 254 40 258 50
rect 262 46 266 60
rect 297 53 300 90
rect 323 77 368 80
rect 319 70 323 77
rect 337 70 341 77
rect 287 49 288 53
rect 293 50 300 53
rect 262 43 284 46
rect 281 40 307 43
rect 254 37 278 40
rect 328 43 332 50
rect 312 39 332 43
rect 340 39 356 43
rect 274 30 278 37
rect 319 30 323 39
rect 330 31 350 35
rect 267 26 279 30
rect 41 15 51 19
rect 78 15 91 19
rect 41 1 44 15
rect 78 10 82 15
rect 144 12 149 14
rect 217 18 247 22
rect 71 6 82 10
rect 41 -3 51 1
rect 78 -32 82 -2
rect 86 -6 90 8
rect 128 8 133 12
rect 144 8 162 12
rect 128 7 129 8
rect 126 1 129 7
rect 144 3 148 8
rect 111 -3 129 1
rect 143 -1 148 3
rect 126 -6 129 -3
rect 126 -10 133 -6
rect 88 -18 138 -15
rect 88 -38 91 -18
rect 99 -26 101 -22
rect 105 -26 113 -22
rect 135 -23 138 -18
rect 127 -27 131 -26
rect 135 -28 136 -23
rect 144 -24 147 -9
rect 151 -15 155 1
rect 217 -6 220 18
rect 274 12 278 19
rect 289 18 303 22
rect 300 12 303 18
rect 267 8 285 12
rect 296 8 303 12
rect 202 -10 227 -6
rect 144 -27 153 -24
rect 100 -38 104 -37
rect 34 -43 47 -40
rect 88 -42 104 -38
rect -165 -63 -140 -59
rect -273 -70 -260 -67
rect -273 -71 -268 -70
rect -291 -75 -268 -74
rect -263 -75 -260 -70
rect -233 -71 -223 -67
rect -187 -71 -175 -67
rect -291 -77 -260 -75
rect -309 -94 -302 -90
rect -291 -91 -287 -77
rect -180 -80 -176 -71
rect -143 -76 -140 -63
rect -17 -51 -11 -48
rect -17 -76 -14 -51
rect -6 -51 27 -48
rect 9 -55 13 -51
rect 27 -55 31 -51
rect 18 -66 22 -65
rect -309 -108 -306 -94
rect -284 -83 -176 -80
rect -152 -79 -14 -76
rect -9 -69 10 -66
rect -9 -77 -6 -69
rect 6 -70 10 -69
rect 18 -70 41 -66
rect 3 -77 20 -73
rect -292 -103 -287 -99
rect -291 -108 -287 -103
rect -284 -101 -280 -83
rect -233 -94 -226 -90
rect -218 -94 -191 -91
rect -309 -112 -302 -108
rect -291 -112 -273 -108
rect -309 -118 -306 -112
rect -309 -122 -295 -118
rect -284 -119 -280 -112
rect -226 -117 -223 -94
rect -309 -149 -306 -122
rect -253 -122 -226 -118
rect -285 -130 -273 -126
rect -284 -133 -280 -130
rect -218 -136 -215 -94
rect -207 -102 -206 -98
rect -195 -99 -191 -94
rect -168 -98 -164 -91
rect -152 -98 -148 -79
rect -141 -99 -137 -91
rect -102 -95 -91 -92
rect -47 -94 -20 -91
rect -102 -98 -99 -95
rect -109 -102 -99 -98
rect -196 -110 -184 -106
rect -142 -110 -129 -106
rect -196 -111 -191 -110
rect -211 -124 -207 -116
rect -196 -117 -191 -116
rect -104 -111 -101 -102
rect -47 -103 -43 -94
rect -54 -107 -42 -103
rect -31 -104 -27 -102
rect -122 -114 -101 -111
rect -196 -121 -184 -117
rect -157 -118 -153 -116
rect -122 -118 -119 -114
rect -85 -116 -81 -114
rect -54 -115 -42 -111
rect -139 -121 -119 -118
rect -211 -130 -207 -128
rect -196 -129 -184 -125
rect -195 -138 -191 -129
rect -215 -141 -191 -138
rect -139 -130 -136 -121
rect -47 -116 -42 -115
rect -31 -116 -27 -108
rect -47 -122 -42 -121
rect -109 -126 -96 -122
rect -54 -126 -42 -122
rect -139 -134 -129 -130
rect -139 -141 -136 -134
rect -101 -141 -97 -133
rect -90 -149 -86 -134
rect -74 -141 -70 -134
rect -47 -138 -43 -133
rect -32 -134 -31 -130
rect -23 -138 -20 -94
rect -47 -141 -25 -138
rect -17 -149 -14 -79
rect 27 -84 31 -70
rect 38 -92 41 -70
rect 44 -84 47 -43
rect 100 -49 104 -42
rect 108 -42 113 -37
rect 118 -42 123 -37
rect 135 -38 138 -28
rect 130 -42 138 -38
rect 108 -49 112 -42
rect 119 -49 123 -42
rect 52 -59 73 -56
rect 52 -63 56 -59
rect 44 -88 63 -84
rect 70 -92 74 -83
rect 78 -81 82 -56
rect 131 -69 138 -65
rect 111 -80 113 -76
rect 131 -85 147 -81
rect 86 -92 90 -91
rect 38 -96 53 -92
rect 61 -96 79 -92
rect 86 -96 102 -92
rect 61 -103 65 -96
rect 86 -103 90 -96
rect 9 -133 13 -124
rect 52 -130 56 -123
rect 70 -130 74 -123
rect 78 -130 82 -123
rect 52 -133 77 -130
rect -309 -152 -14 -149
rect 9 -139 13 -138
rect 68 -139 71 -133
rect 9 -142 86 -139
rect 9 -149 13 -142
rect -312 -158 -2 -155
rect -5 -197 -2 -158
rect 37 -169 41 -142
rect 68 -149 72 -142
rect 86 -149 90 -142
rect 77 -176 81 -169
rect 56 -180 69 -176
rect 77 -180 96 -176
rect 27 -196 31 -189
rect 45 -196 49 -189
rect 56 -196 59 -180
rect -5 -200 20 -197
rect 27 -200 38 -196
rect 45 -200 59 -196
rect 62 -188 79 -184
rect 27 -203 31 -200
rect 3 -207 10 -203
rect 18 -207 31 -203
rect 45 -201 49 -200
rect 62 -203 65 -188
rect 86 -189 90 -180
rect 59 -206 65 -203
rect 93 -203 96 -180
rect 99 -196 102 -96
rect 119 -104 123 -91
rect 130 -96 136 -92
rect 144 -118 147 -85
rect 127 -131 131 -124
rect 150 -127 153 -27
rect 176 -106 180 -10
rect 275 -21 278 1
rect 281 3 285 8
rect 300 6 303 8
rect 281 -1 286 3
rect 300 2 314 6
rect 337 6 341 10
rect 319 3 341 6
rect 300 -6 303 2
rect 319 -1 323 3
rect 337 -1 341 3
rect 347 -2 350 31
rect 281 -13 285 -9
rect 296 -10 303 -6
rect 328 -12 332 -11
rect 347 -12 350 -7
rect 281 -16 306 -13
rect 311 -16 332 -12
rect 340 -16 350 -12
rect 353 25 356 39
rect 353 20 357 25
rect 157 -109 180 -106
rect 127 -139 131 -136
rect 157 -139 160 -109
rect 176 -116 180 -109
rect 222 -24 278 -21
rect 109 -142 160 -139
rect 109 -149 113 -142
rect 137 -169 141 -142
rect 170 -148 177 -144
rect 184 -149 188 -136
rect 162 -159 176 -155
rect 194 -164 196 -160
rect 169 -175 176 -171
rect 127 -196 131 -189
rect 145 -196 149 -189
rect 99 -200 120 -196
rect 127 -200 138 -196
rect 145 -199 166 -196
rect 184 -198 188 -191
rect 195 -198 199 -191
rect 145 -200 177 -199
rect 127 -203 131 -200
rect 3 -228 6 -207
rect 18 -208 22 -207
rect 9 -222 13 -218
rect 27 -222 31 -218
rect 37 -220 41 -211
rect 9 -225 36 -222
rect 2 -241 6 -233
rect 21 -241 24 -225
rect 59 -226 62 -206
rect 93 -207 110 -203
rect 118 -207 131 -203
rect 145 -201 149 -200
rect 163 -202 177 -200
rect 68 -220 72 -209
rect 118 -208 122 -207
rect 109 -222 113 -218
rect 127 -222 131 -218
rect 137 -222 141 -211
rect 72 -225 157 -222
rect 169 -222 172 -202
rect 184 -203 189 -198
rect 194 -203 199 -198
rect 203 -198 207 -191
rect 203 -202 219 -198
rect 203 -203 207 -202
rect 176 -214 180 -213
rect 194 -218 202 -214
rect 206 -218 208 -214
rect 216 -222 219 -202
rect 169 -225 219 -222
rect 58 -228 62 -226
rect 222 -228 225 -24
rect 319 -30 323 -16
rect 353 -19 356 20
rect 330 -23 356 -19
rect 365 -30 368 77
rect 341 -34 368 -30
rect 58 -231 225 -228
rect 58 -241 61 -231
rect -12 -245 6 -241
rect 17 -245 24 -241
rect 48 -245 61 -241
rect 88 -245 95 -241
rect -16 -288 -12 -263
rect -5 -275 -1 -252
rect 2 -250 6 -245
rect 2 -254 7 -250
rect 21 -259 24 -245
rect 2 -269 6 -262
rect 17 -263 28 -259
rect 2 -272 11 -269
rect 49 -269 53 -252
rect 58 -250 61 -245
rect 58 -254 68 -250
rect 16 -272 53 -269
rect 95 -259 98 -245
rect 57 -275 61 -262
rect 88 -263 98 -259
rect -5 -278 61 -275
rect 34 -280 39 -278
rect 95 -288 98 -263
rect -16 -291 98 -288
<< m2contact >>
rect 20 267 25 272
rect 116 259 121 264
rect 29 230 34 235
rect -95 144 -90 149
rect -166 124 -161 129
rect -95 125 -90 130
rect -95 111 -90 116
rect 84 184 89 189
rect 30 168 35 173
rect -15 135 -10 140
rect -138 100 -133 105
rect -95 79 -90 84
rect -166 59 -161 64
rect -150 60 -145 65
rect -95 60 -90 65
rect -317 12 -312 17
rect -356 2 -351 7
rect -95 46 -90 51
rect -138 35 -133 40
rect -111 39 -106 44
rect -56 57 -51 62
rect 71 145 76 150
rect 95 144 100 149
rect 118 184 123 189
rect 95 117 100 122
rect 51 74 56 79
rect 70 74 75 79
rect 84 74 89 79
rect 150 82 155 87
rect 254 72 259 77
rect -32 29 -27 34
rect -161 16 -156 21
rect -152 13 -147 18
rect -136 -13 -131 -8
rect 44 53 49 58
rect -76 -14 -71 -9
rect -57 -14 -52 -9
rect -43 -14 -38 -9
rect 78 50 84 56
rect -318 -44 -313 -39
rect -143 -37 -138 -32
rect -5 -38 0 -33
rect 126 24 131 29
rect 208 44 213 49
rect 318 77 323 82
rect 307 39 312 44
rect 144 14 149 19
rect 86 -11 92 -6
rect 76 -37 82 -32
rect 94 -26 99 -21
rect 113 -26 118 -21
rect 127 -26 132 -21
rect 136 -28 141 -23
rect 150 -20 155 -15
rect -268 -75 -263 -70
rect 27 -51 32 -46
rect -169 -91 -164 -86
rect -285 -138 -280 -133
rect -212 -102 -207 -97
rect -91 -95 -86 -90
rect -212 -116 -207 -111
rect -157 -116 -152 -111
rect -141 -115 -136 -110
rect -31 -102 -26 -97
rect -211 -135 -206 -130
rect -221 -142 -215 -136
rect -102 -122 -97 -117
rect -86 -121 -81 -116
rect -31 -121 -26 -116
rect -101 -146 -96 -141
rect -31 -134 -26 -129
rect -74 -146 -69 -141
rect -11 -82 -6 -77
rect 73 -60 78 -55
rect 138 -69 143 -64
rect 8 -138 13 -133
rect 77 -135 82 -130
rect -317 -158 -312 -153
rect 114 -97 119 -92
rect 142 -123 147 -118
rect 345 -7 350 -2
rect 306 -17 311 -12
rect 126 -136 132 -131
rect 149 -132 154 -127
rect 188 -148 193 -143
rect 157 -160 162 -155
rect 164 -176 169 -171
rect 36 -225 41 -220
rect 67 -225 72 -220
rect 157 -225 162 -220
rect 175 -219 180 -214
rect 189 -219 194 -214
rect 208 -219 213 -214
rect 11 -272 16 -267
<< metal2 >>
rect 21 284 107 287
rect 21 272 24 284
rect -84 233 -58 234
rect -84 231 29 233
rect -165 144 -95 147
rect -165 129 -162 144
rect -148 105 -145 125
rect -95 116 -91 125
rect -160 102 -138 105
rect -165 79 -95 82
rect -165 64 -162 79
rect -148 40 -145 60
rect -95 51 -91 60
rect -160 37 -138 40
rect -111 31 -107 39
rect -168 29 -107 31
rect -371 28 -107 29
rect -371 26 -165 28
rect -371 6 -368 26
rect -84 24 -81 231
rect -63 230 29 231
rect 30 173 34 230
rect 89 184 90 189
rect 53 146 71 149
rect -10 137 35 140
rect -39 96 13 99
rect -150 21 -81 24
rect -74 58 -56 61
rect -316 17 -161 20
rect -150 18 -147 21
rect -317 9 -306 12
rect -371 3 -356 6
rect -316 -153 -313 -44
rect -309 -79 -306 9
rect -74 -9 -71 58
rect -32 44 -29 56
rect 9 54 13 96
rect 32 58 35 137
rect 53 79 56 146
rect 95 132 98 144
rect 75 129 98 132
rect 95 122 98 129
rect 104 122 107 284
rect 118 189 121 259
rect 117 184 118 189
rect 100 119 107 122
rect 119 82 150 85
rect 75 75 84 79
rect 32 55 44 58
rect 119 56 122 82
rect 300 77 318 80
rect 84 53 122 56
rect 213 45 280 48
rect -52 41 -29 44
rect -32 34 -29 41
rect -18 40 129 43
rect -135 -32 -132 -13
rect -52 -13 -43 -9
rect -138 -35 -132 -32
rect -18 -72 -15 40
rect 126 29 129 40
rect 277 42 280 45
rect 300 42 303 77
rect 277 39 303 42
rect 116 16 144 19
rect 116 -6 119 16
rect 92 -9 119 -6
rect 350 -6 365 -3
rect 155 -20 310 -17
rect 118 -26 127 -22
rect 0 -37 76 -34
rect 32 -51 76 -48
rect 73 -55 76 -51
rect -263 -75 -15 -72
rect -309 -82 -11 -79
rect -164 -91 -142 -88
rect -91 -89 -10 -86
rect -91 -90 -86 -89
rect -211 -111 -207 -102
rect -157 -111 -154 -91
rect -101 -102 -31 -99
rect -140 -130 -137 -115
rect -101 -117 -98 -102
rect -206 -133 -137 -130
rect -280 -138 -221 -137
rect -285 -140 -221 -138
rect -84 -141 -81 -121
rect -31 -129 -27 -121
rect -13 -133 -10 -89
rect 74 -120 77 -60
rect 96 -93 99 -26
rect 362 -24 365 -6
rect 141 -27 365 -24
rect 138 -76 141 -69
rect 118 -79 141 -76
rect 138 -91 141 -79
rect 96 -96 114 -93
rect 74 -123 142 -120
rect 147 -122 161 -119
rect -13 -136 8 -133
rect 82 -131 111 -130
rect 82 -133 126 -131
rect 99 -134 126 -133
rect -96 -144 -74 -141
rect -99 -150 -96 -146
rect -99 -153 -8 -150
rect -11 -284 -8 -153
rect 41 -225 67 -222
rect 150 -230 153 -132
rect 158 -155 161 -122
rect 193 -147 211 -144
rect 157 -220 160 -160
rect 166 -161 169 -149
rect 166 -164 189 -161
rect 166 -171 169 -164
rect 208 -214 211 -147
rect 180 -218 189 -214
rect 7 -233 153 -230
rect 12 -284 15 -272
rect -11 -287 15 -284
<< m123contact >>
rect -7 278 -2 283
rect -64 241 -59 246
rect 11 239 16 244
rect -150 125 -145 130
rect -111 125 -106 130
rect -165 100 -160 105
rect -111 60 -106 65
rect -165 35 -160 40
rect 89 231 94 236
rect -72 222 -67 227
rect -23 153 -18 158
rect -44 96 -39 101
rect -369 -25 -362 -19
rect -330 -82 -325 -77
rect -32 56 -27 61
rect -57 41 -52 46
rect 70 129 75 134
rect 215 145 220 150
rect 70 90 75 95
rect 92 90 97 95
rect 123 93 128 98
rect 208 93 213 98
rect -25 47 -20 52
rect 8 49 14 54
rect 208 59 213 64
rect 288 48 293 53
rect -57 2 -52 7
rect -302 -22 -297 -17
rect -155 -22 -150 -17
rect -128 -39 -123 -34
rect -302 -53 -297 -48
rect -226 -61 -214 -56
rect 40 26 45 31
rect 133 33 138 38
rect 357 20 362 25
rect 123 7 128 12
rect 314 2 319 7
rect -11 -53 -6 -48
rect -2 -77 3 -72
rect -226 -94 -221 -89
rect -142 -91 -137 -86
rect -196 -116 -191 -111
rect -226 -122 -221 -117
rect -47 -121 -42 -116
rect 113 -42 118 -37
rect 113 -81 118 -76
rect 136 -96 141 -91
rect -141 -146 -136 -141
rect -25 -143 -20 -138
rect 86 -142 92 -137
rect 2 -233 7 -228
rect 165 -149 170 -144
rect 189 -164 194 -159
rect 189 -203 194 -198
rect 95 -245 100 -240
rect 34 -285 39 -280
<< metal3 >>
rect -2 280 103 283
rect -73 241 -64 244
rect -73 227 -70 241
rect 11 236 16 239
rect -21 233 89 236
rect -73 224 -72 227
rect -116 153 -113 159
rect -116 150 -108 153
rect -111 130 -108 150
rect -163 88 -160 100
rect -70 99 -67 222
rect -21 158 -18 233
rect -70 96 -44 99
rect 100 95 103 280
rect 211 145 215 148
rect 210 98 213 145
rect 24 92 70 95
rect -163 85 -108 88
rect -111 65 -108 85
rect 24 61 27 92
rect 97 92 103 95
rect -27 58 27 61
rect -20 47 -8 50
rect 14 49 44 52
rect -165 28 -162 35
rect -369 25 -162 28
rect -369 -19 -366 25
rect -80 7 -77 12
rect -80 4 -57 7
rect -150 -22 -125 -19
rect -302 -48 -299 -22
rect -128 -34 -125 -22
rect -11 -48 -8 47
rect 41 31 44 49
rect 123 36 126 93
rect 208 64 211 93
rect 123 33 133 36
rect 288 36 291 48
rect 212 33 318 36
rect 123 23 126 33
rect 212 23 215 33
rect 123 20 215 23
rect 123 12 126 20
rect 315 7 318 33
rect 362 20 363 25
rect 360 -18 363 20
rect 157 -21 363 -18
rect 90 -42 113 -39
rect -222 -76 -219 -61
rect -225 -77 -219 -76
rect -325 -79 -219 -77
rect -325 -80 -222 -79
rect -225 -89 -222 -80
rect -95 -86 -44 -83
rect -95 -88 -92 -86
rect -137 -91 -92 -88
rect -225 -143 -222 -122
rect -194 -136 -191 -116
rect -47 -116 -44 -86
rect -194 -139 -186 -136
rect -225 -146 -141 -143
rect -23 -148 -20 -143
rect -23 -151 -6 -148
rect -9 -284 -6 -151
rect -1 -231 2 -77
rect 90 -130 93 -42
rect 157 -91 160 -21
rect 141 -94 160 -91
rect 90 -133 106 -130
rect 103 -137 106 -133
rect 92 -142 99 -139
rect 103 -140 168 -137
rect 96 -240 99 -142
rect 165 -144 168 -140
rect 214 -198 217 -193
rect 194 -201 217 -198
rect -9 -285 34 -284
rect -9 -287 38 -285
<< m234contact >>
rect 90 184 95 189
rect 112 184 117 189
rect 206 145 211 150
<< metal4 >>
rect 95 184 112 187
rect 112 148 115 184
rect 112 145 206 148
<< labels >>
rlabel metal3 91 -53 91 -53 1 node31
rlabel metal3 -53 -85 -49 -84 1 node21
rlabel metal3 -122 86 -118 87 1 node11
rlabel metal3 39 93 40 94 1 node01
rlabel metal1 79 21 81 26 1 Pout_bar
rlabel metal1 146 11 146 11 1 node34
rlabel metal1 172 74 172 74 1 node35
rlabel metal1 256 69 256 69 1 node33
rlabel metal1 276 30 276 30 1 node32
rlabel metal2 357 -5 359 -4 1 B3
rlabel metal1 354 20 355 23 1 A3
rlabel metal1 164 -198 164 -198 1 C3
rlabel metal1 -63 183 -63 183 1 C1
rlabel metal1 95 -95 95 -95 1 node25
rlabel metal1 92 -179 92 -179 1 node23
rlabel metal1 34 -69 34 -69 1 node24
rlabel metal1 52 -199 52 -199 1 node22
rlabel metal2 13 -281 14 -279 1 B2
rlabel metal1 -282 -131 -282 -131 1 C2
rlabel metal1 -262 -69 -262 -69 1 node13
rlabel metal1 -179 -76 -179 -76 1 node15
rlabel metal1 -152 -16 -152 -16 1 node14
rlabel metal1 -283 -35 -283 -35 1 node12
rlabel metal1 -361 -23 -360 -21 1 A1
rlabel metal1 -28 171 -28 171 1 node02
rlabel metal1 140 199 146 202 1 gnd
rlabel metal1 140 185 146 188 1 vdd
rlabel metal1 -5 284 -4 286 1 A0
rlabel metal2 22 284 23 285 1 B0
rlabel metal3 -115 153 -114 158 1 S1
rlabel metal1 35 -278 38 -276 1 A2
rlabel metal3 215 -197 216 -194 1 S3
rlabel metal3 -190 -138 -187 -137 1 S2
rlabel metal3 -79 8 -78 11 1 S0
rlabel metal1 255 158 257 160 1 Cout
rlabel metal1 151 137 153 139 1 node36
rlabel metal1 275 114 277 117 1 Gout_bar
rlabel metal1 315 40 317 42 1 G3_bar
rlabel metal1 315 -15 317 -13 1 P3_bar
rlabel metal1 3 -239 5 -237 1 P2_bar
rlabel metal1 58 -239 60 -237 1 G2_bar
rlabel metal1 -323 -42 -321 -40 1 G1_bar
rlabel metal1 -323 13 -321 15 1 P1_bar
rlabel metal2 -366 4 -363 5 1 B1
rlabel metal1 31 237 33 239 1 P0_bar
rlabel metal1 -24 237 -22 239 1 G0_bar
rlabel metal1 24 -1 26 1 1 C0_bar
rlabel metal1 -1 -1 1 1 1 C0
<< end >>
