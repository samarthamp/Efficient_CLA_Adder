* SPICE3 file created from /home/mpsamartha/Ubuntu_Backed/Project/Magic/pg_layout.ext - technology: scmos

.option scale=0.09u

M1000 G_bar A vdd w_n69_n66# pfet w=20 l=2
+  ad=160 pd=56 as=400 ps=190
M1001 vdd B G_bar w_n69_n66# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 P_bar B gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=200 ps=110
M1003 a_n56_n20# A gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1004 a_n56_40# B vdd w_n69_34# pfet w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1005 gnd A P_bar Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 G_bar B a_n56_n20# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1007 P_bar A a_n56_40# w_n69_34# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
C0 w_n69_34# P_bar 0.02fF
C1 A B 1.25fF
C2 w_n69_34# B 0.06fF
C3 P_bar gnd 0.02fF
C4 A G_bar 0.04fF
C5 w_n69_n66# vdd 0.05fF
C6 gnd B 0.15fF
C7 P_bar B 0.04fF
C8 w_n69_n66# A 0.07fF
C9 w_n69_34# vdd 0.02fF
C10 G_bar B 0.19fF
C11 w_n69_34# A 0.06fF
C12 w_n69_n66# B 0.07fF
C13 A P_bar 0.21fF
C14 w_n69_n66# G_bar 0.02fF
C15 vdd Gnd 0.08fF
C16 G_bar Gnd 0.09fF
C17 gnd Gnd 0.11fF
C18 P_bar Gnd 0.05fF
C19 A Gnd 0.34fF
C20 B Gnd 0.46fF
C21 w_n69_n66# Gnd 1.03fF
C22 w_n69_34# Gnd 1.78fF
