* SPICE3 file created from nand_layout.ext - technology: scmos

.include TSMC_180nm.txt
.param vdd=1.8
.param LAMBDA=0.09u
.global vdd gnd
.option scale=0.09u

M1000 out b a_13_n34# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=160 ps=56
M1001 out a vdd w_0_0# CMOSP w=20 l=2
+  ad=160 pd=56 as=200 ps=100
M1002 a_13_n34# a gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1003 vdd b out w_0_0# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 b a 0.21fF
C1 w_0_0# out 0.02fF
C2 a out 0.04fF
C3 w_0_0# a 0.07fF
C4 b out 0.19fF
C5 w_0_0# vdd 0.05fF
C6 b w_0_0# 0.07fF

Vdd vdd gnd dc 1.8
* trise = tfall = 5% of T_on
Va  a  gnd pulse 1.8 0 10ns 100ps   100ps   20ns 40ns
Vb  b  gnd pulse 1.8 0 10ns 100ps   100ps   40ns 80ns
* .ic v(out) = 0
.tran 1ps 200ns 1ps
* CL out gnd 50f

* clk - out propagation delay
.measure tran t_rise TRIG V(a) VAL='0.9' FALL=1 TARG V(out) VAL='0.9' RISE=1
.measure tran t_fall TRIG V(a) VAL='0.9' RISE=2 TARG V(out) VAL='0.9' FALL=1
.measure tran prop_delay param ='(t_rise + t_fall)/2'

* 20lambda: 304p, 245p, 275p
* saturates around 90p

.control
set hcopypscolor = 1
set color0 = white
set color1 = black

run
set curplottitle= "M P Samartha-2023102038"
plot a+4, b+2, out
.endc



