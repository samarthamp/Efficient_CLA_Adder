* SPICE3 file created from xor.ext - technology: scmos

.include TSMC_180nm.txt
.param vdd=1.8
.param LAMBDA=0.09u
.global vdd gnd
.option scale=0.09u

M1000 a_39_n44# a_bar out Gnd CMOSN w=30 l=2
+  ad=240 pd=76 as=420 ps=88
M1001 a_13_n44# a gnd Gnd CMOSN w=30 l=2
+  ad=240 pd=76 as=400 ps=200
M1002 a_13_6# a vdd w_0_0# CMOSP w=40 l=2
+  ad=720 pd=276 as=600 ps=280
M1003 b_bar b vdd w_n39_n58# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1004 out a_bar a_13_6# w_0_0# CMOSP w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1005 vdd b a_13_6# w_0_0# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 a_13_6# b_bar out w_0_0# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_bar a gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1008 gnd b_bar a_39_n44# Gnd CMOSN w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 b_bar b gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1010 out b a_13_n44# Gnd CMOSN w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 a_bar a vdd w_n39_21# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 a_13_6# b 0.12fF
C1 a_13_6# a_bar 0.13fF
C2 b gnd 0.14fF
C3 vdd b 0.07fF
C4 a_bar vdd 0.06fF
C5 w_0_0# b_bar 0.06fF
C6 w_n39_n58# b 0.07fF
C7 w_0_0# a 0.06fF
C8 w_n39_21# vdd 0.02fF
C9 out b_bar 0.06fF
C10 a_13_6# vdd 0.14fF
C11 out w_0_0# 0.02fF
C12 b b_bar 0.10fF
C13 a b 0.13fF
C14 w_n39_n58# vdd 0.02fF
C15 a_bar a 0.05fF
C16 w_0_0# b 0.06fF
C17 w_n39_21# a 0.07fF
C18 w_0_0# a_bar 0.08fF
C19 out b 0.04fF
C20 a_13_6# a 0.04fF
C21 out a_bar 0.06fF
C22 a_13_6# w_0_0# 0.09fF
C23 a_13_6# out 0.20fF
C24 b_bar gnd 0.28fF
C25 a gnd 0.13fF
C26 w_n39_n58# b_bar 0.02fF
C27 a vdd 0.07fF
C28 w_0_0# vdd 0.05fF
C29 w_n39_21# a_bar 0.02fF
C30 out Gnd 0.12fF
C31 a_13_6# Gnd 0.06fF
C32 gnd Gnd 0.17fF
C33 b_bar Gnd 1.38fF
C34 b Gnd 0.93fF
C35 vdd Gnd 0.61fF
C36 a Gnd 0.97fF
C37 a_bar Gnd 0.29fF
C38 w_n39_n58# Gnd 0.77fF
C39 w_0_0# Gnd 0.99fF
C40 w_n39_21# Gnd 0.77fF

Vdd vdd gnd dc 1.8
* trise = tfall = 5% of T_on
Va  a  gnd pulse 1.8 0 5n 100ps  100ps  10ns 20ns
Vb  b  gnd pulse 1.8 0 0  100ps  100ps  20ns 40ns
* .ic v(out) = 0
.tran 100ps 200ns 1ps
* CL out gnd 50f

* clk - out propagation delay
.measure tran t_rise TRIG V(a) VAL='0.9' FALL=1 TARG V(out) VAL='0.9' RISE=1
.measure tran t_fall TRIG V(a) VAL='0.9' RISE=2 TARG V(out) VAL='0.9' FALL=1
.measure tran prop_delay param ='(t_rise + t_fall)/2'

* 20lambda: 304p, 245p, 275p
* saturates around 90p

.control
set hcopypscolor = 1
set color0 = white
set color1 = black

run
set curplottitle= "M P Samartha-2023102038"
plot a+4, b+2, out
.endc





